VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/"  ;

SITE TSM130NMMETROSITE
    SYMMETRY Y  ;
    CLASS core  ;
    SIZE 0.410 BY 2.870 ;
END TSM130NMMETROSITE

MACRO ADDFHX1MTH
    CLASS CORE ;
    FOREIGN ADDFHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.220 0.730 11.380 2.140 ;
        RECT  11.090 0.730 11.220 0.990 ;
        RECT  11.090 1.700 11.220 2.140 ;
        END
        AntennaDiffArea 0.333 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.350 0.705 10.560 1.880 ;
        RECT  10.145 0.705 10.350 0.965 ;
        RECT  10.060 1.720 10.350 1.880 ;
        END
        AntennaDiffArea 0.329 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.120 0.880 9.400 1.615 ;
        END
        AntennaGateArea 0.1534 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.290 5.325 1.765 ;
        END
        AntennaGateArea 0.5876 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.090 0.485 1.580 ;
        END
        AntennaGateArea 0.26 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.065 -0.130 11.480 0.130 ;
        RECT  10.465 -0.130 11.065 0.300 ;
        RECT  1.675 -0.130 10.465 0.130 ;
        RECT  0.735 -0.130 1.675 0.250 ;
        RECT  0.000 -0.130 0.735 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.200 2.740 11.480 3.000 ;
        RECT  10.600 2.555 11.200 3.000 ;
        RECT  5.525 2.740 10.600 3.000 ;
        RECT  5.265 2.285 5.525 3.000 ;
        RECT  1.500 2.740 5.265 3.000 ;
        RECT  0.900 2.265 1.500 3.000 ;
        RECT  0.000 2.740 0.900 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.900 1.230 11.035 1.490 ;
        RECT  10.740 1.230 10.900 2.220 ;
        RECT  8.215 2.060 10.740 2.220 ;
        RECT  6.645 2.400 10.395 2.560 ;
        RECT  9.810 0.540 9.895 0.945 ;
        RECT  9.635 0.540 9.810 1.880 ;
        RECT  9.390 0.540 9.635 0.700 ;
        RECT  9.550 1.720 9.635 1.880 ;
        RECT  9.230 0.310 9.390 0.700 ;
        RECT  7.875 0.310 9.230 0.470 ;
        RECT  8.740 0.725 8.900 1.880 ;
        RECT  8.395 1.720 8.740 1.880 ;
        RECT  8.215 0.735 8.440 0.895 ;
        RECT  8.055 0.735 8.215 2.220 ;
        RECT  7.885 1.960 8.055 2.220 ;
        RECT  7.715 0.310 7.875 0.945 ;
        RECT  7.705 0.785 7.715 0.945 ;
        RECT  7.545 0.785 7.705 1.935 ;
        RECT  7.085 1.775 7.545 1.935 ;
        RECT  7.025 0.310 7.510 0.470 ;
        RECT  7.205 0.685 7.365 1.595 ;
        RECT  6.645 1.435 7.205 1.595 ;
        RECT  6.825 1.775 7.085 2.155 ;
        RECT  6.865 0.310 7.025 1.255 ;
        RECT  3.885 0.310 6.865 0.470 ;
        RECT  6.245 1.095 6.865 1.255 ;
        RECT  6.525 0.655 6.685 0.915 ;
        RECT  6.485 1.435 6.645 2.560 ;
        RECT  5.865 0.685 6.525 0.845 ;
        RECT  6.285 2.165 6.485 2.425 ;
        RECT  6.085 1.095 6.245 1.975 ;
        RECT  5.865 2.165 6.035 2.425 ;
        RECT  5.705 0.685 5.865 2.425 ;
        RECT  5.515 0.685 5.705 0.845 ;
        RECT  5.015 1.945 5.705 2.105 ;
        RECT  5.165 0.650 5.325 1.035 ;
        RECT  4.225 0.650 5.165 0.810 ;
        RECT  4.795 1.945 5.015 2.345 ;
        RECT  4.635 1.625 4.795 2.345 ;
        RECT  4.455 0.990 4.695 1.385 ;
        RECT  4.435 0.990 4.455 2.560 ;
        RECT  4.295 1.225 4.435 2.560 ;
        RECT  2.275 2.400 4.295 2.560 ;
        RECT  4.115 0.650 4.225 1.045 ;
        RECT  4.065 0.650 4.115 2.220 ;
        RECT  3.955 0.885 4.065 2.220 ;
        RECT  2.785 2.060 3.955 2.220 ;
        RECT  3.775 0.310 3.885 0.705 ;
        RECT  3.615 0.310 3.775 1.880 ;
        RECT  3.515 1.720 3.615 1.880 ;
        RECT  3.165 0.430 3.325 1.880 ;
        RECT  0.890 0.430 3.165 0.590 ;
        RECT  3.005 1.720 3.165 1.880 ;
        RECT  2.625 0.800 2.785 2.220 ;
        RECT  2.525 0.800 2.625 0.960 ;
        RECT  2.495 1.880 2.625 2.220 ;
        RECT  2.115 0.795 2.275 2.560 ;
        RECT  2.015 0.795 2.115 0.955 ;
        RECT  1.985 1.825 2.115 2.560 ;
        RECT  1.365 1.285 1.900 1.545 ;
        RECT  1.205 0.815 1.365 1.945 ;
        RECT  1.105 0.815 1.205 0.975 ;
        RECT  1.075 1.685 1.205 1.945 ;
        RECT  0.730 0.430 0.890 2.005 ;
        RECT  0.125 0.645 0.730 0.905 ;
        RECT  0.385 1.760 0.730 2.005 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END ADDFHX1MTH

MACRO ADDFHX2MTH
    CLASS CORE ;
    FOREIGN ADDFHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.450 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.315 1.290 18.350 1.580 ;
        RECT  18.300 0.420 18.315 1.580 ;
        RECT  18.140 0.420 18.300 2.100 ;
        RECT  18.055 0.420 18.140 1.020 ;
        RECT  17.770 1.940 18.140 2.100 ;
        RECT  17.610 1.940 17.770 2.420 ;
        RECT  17.510 2.160 17.610 2.420 ;
        END
        AntennaDiffArea 0.399 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.135 0.410 17.235 0.670 ;
        RECT  16.975 0.410 17.135 1.170 ;
        RECT  16.910 0.880 16.975 1.170 ;
        RECT  16.675 1.010 16.910 1.170 ;
        RECT  16.515 1.010 16.675 1.760 ;
        RECT  16.305 1.600 16.515 1.760 ;
        END
        AntennaDiffArea 0.492 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.090 0.880 16.300 1.170 ;
        RECT  15.885 1.010 16.090 1.170 ;
        RECT  15.615 1.010 15.885 1.330 ;
        END
        AntennaGateArea 0.2418 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.560 1.450 10.805 1.710 ;
        RECT  10.350 1.290 10.560 1.710 ;
        RECT  10.205 1.450 10.350 1.710 ;
        END
        AntennaGateArea 0.9386 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.230 0.945 1.490 ;
        RECT  0.100 1.230 0.310 1.580 ;
        END
        AntennaGateArea 0.4264 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.775 -0.130 18.450 0.130 ;
        RECT  17.515 -0.130 17.775 0.980 ;
        RECT  16.725 -0.130 17.515 0.130 ;
        RECT  16.465 -0.130 16.725 0.670 ;
        RECT  15.625 -0.130 16.465 0.130 ;
        RECT  15.465 -0.130 15.625 0.300 ;
        RECT  11.345 -0.130 15.465 0.130 ;
        RECT  10.405 -0.130 11.345 0.250 ;
        RECT  2.645 -0.130 10.405 0.130 ;
        RECT  2.045 -0.130 2.645 0.250 ;
        RECT  1.665 -0.130 2.045 0.130 ;
        RECT  1.065 -0.130 1.665 0.250 ;
        RECT  0.385 -0.130 1.065 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.280 2.740 18.450 3.000 ;
        RECT  18.020 2.280 18.280 3.000 ;
        RECT  17.170 2.740 18.020 3.000 ;
        RECT  16.910 2.280 17.170 3.000 ;
        RECT  15.030 2.740 16.910 3.000 ;
        RECT  14.770 2.620 15.030 3.000 ;
        RECT  10.585 2.740 14.770 3.000 ;
        RECT  10.325 2.235 10.585 3.000 ;
        RECT  9.565 2.740 10.325 3.000 ;
        RECT  9.305 2.235 9.565 3.000 ;
        RECT  2.675 2.740 9.305 3.000 ;
        RECT  2.415 2.200 2.675 3.000 ;
        RECT  1.325 2.740 2.415 3.000 ;
        RECT  1.065 2.570 1.325 3.000 ;
        RECT  0.725 2.740 1.065 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.340 1.425 17.940 1.685 ;
        RECT  17.220 1.525 17.340 1.685 ;
        RECT  17.060 1.525 17.220 2.100 ;
        RECT  13.625 1.940 17.060 2.100 ;
        RECT  15.955 0.440 16.215 0.700 ;
        RECT  12.705 2.280 16.195 2.440 ;
        RECT  15.285 0.490 15.955 0.650 ;
        RECT  15.285 1.600 15.645 1.760 ;
        RECT  15.125 0.330 15.285 1.760 ;
        RECT  13.925 0.330 15.125 0.490 ;
        RECT  14.875 1.600 15.125 1.760 ;
        RECT  14.845 0.680 14.945 0.890 ;
        RECT  14.610 1.450 14.875 1.760 ;
        RECT  14.685 0.680 14.845 1.270 ;
        RECT  14.330 1.110 14.685 1.270 ;
        RECT  14.175 0.680 14.435 0.930 ;
        RECT  14.170 1.110 14.330 1.760 ;
        RECT  13.625 0.770 14.175 0.930 ;
        RECT  14.070 1.550 14.170 1.760 ;
        RECT  13.665 0.330 13.925 0.575 ;
        RECT  12.915 0.330 13.665 0.490 ;
        RECT  13.465 0.770 13.625 2.100 ;
        RECT  13.355 0.770 13.465 0.930 ;
        RECT  13.095 0.670 13.355 0.930 ;
        RECT  13.115 1.820 13.215 2.080 ;
        RECT  12.955 1.360 13.115 2.080 ;
        RECT  12.915 1.360 12.955 1.520 ;
        RECT  12.755 0.330 12.915 1.520 ;
        RECT  12.525 0.500 12.755 0.760 ;
        RECT  12.575 1.900 12.705 2.560 ;
        RECT  12.415 1.130 12.575 2.560 ;
        RECT  12.275 1.130 12.415 1.290 ;
        RECT  11.555 2.400 12.415 2.560 ;
        RECT  12.115 0.500 12.275 1.290 ;
        RECT  12.075 1.470 12.235 1.880 ;
        RECT  12.065 0.500 12.115 0.760 ;
        RECT  11.895 2.060 12.115 2.220 ;
        RECT  11.885 1.470 12.075 1.630 ;
        RECT  11.735 1.810 11.895 2.220 ;
        RECT  11.725 0.310 11.885 1.630 ;
        RECT  11.205 1.810 11.735 1.970 ;
        RECT  11.625 0.310 11.725 0.590 ;
        RECT  9.725 0.430 11.625 0.590 ;
        RECT  11.395 2.150 11.555 2.560 ;
        RECT  11.385 0.770 11.545 1.580 ;
        RECT  8.155 0.770 11.385 0.930 ;
        RECT  11.095 1.110 11.205 2.055 ;
        RECT  11.045 1.110 11.095 2.375 ;
        RECT  10.945 1.110 11.045 1.270 ;
        RECT  10.835 1.895 11.045 2.375 ;
        RECT  10.075 1.895 10.835 2.055 ;
        RECT  10.025 1.110 10.125 1.270 ;
        RECT  10.025 1.895 10.075 2.495 ;
        RECT  9.865 1.110 10.025 2.495 ;
        RECT  9.815 1.895 9.865 2.495 ;
        RECT  9.055 1.895 9.815 2.055 ;
        RECT  9.465 0.385 9.725 0.590 ;
        RECT  7.815 0.385 9.465 0.545 ;
        RECT  8.495 1.110 9.185 1.270 ;
        RECT  8.955 1.895 9.055 2.495 ;
        RECT  8.795 1.450 8.955 2.495 ;
        RECT  8.705 1.450 8.795 1.710 ;
        RECT  8.335 1.110 8.495 2.560 ;
        RECT  4.205 2.400 8.335 2.560 ;
        RECT  7.995 0.770 8.155 2.220 ;
        RECT  5.585 2.060 7.995 2.220 ;
        RECT  7.655 0.385 7.815 1.880 ;
        RECT  7.385 0.385 7.655 0.645 ;
        RECT  6.375 1.720 7.655 1.880 ;
        RECT  7.225 0.385 7.385 0.925 ;
        RECT  6.125 1.380 7.355 1.540 ;
        RECT  6.435 0.765 7.225 0.925 ;
        RECT  6.715 0.310 6.975 0.585 ;
        RECT  5.845 0.310 6.715 0.470 ;
        RECT  6.175 0.650 6.435 0.925 ;
        RECT  5.865 1.380 6.125 1.880 ;
        RECT  5.845 1.380 5.865 1.600 ;
        RECT  5.685 0.310 5.845 1.600 ;
        RECT  4.845 0.310 5.685 0.470 ;
        RECT  5.035 1.440 5.685 1.600 ;
        RECT  5.325 1.835 5.585 2.220 ;
        RECT  4.595 2.060 5.325 2.220 ;
        RECT  5.145 0.685 5.305 1.235 ;
        RECT  3.755 1.075 5.145 1.235 ;
        RECT  4.875 1.440 5.035 1.880 ;
        RECT  4.775 1.720 4.875 1.880 ;
        RECT  4.585 0.310 4.845 0.895 ;
        RECT  4.435 1.880 4.595 2.220 ;
        RECT  2.985 0.310 4.585 0.470 ;
        RECT  3.695 1.880 4.435 2.040 ;
        RECT  3.315 0.650 4.295 0.810 ;
        RECT  3.945 2.220 4.205 2.560 ;
        RECT  3.185 2.330 3.945 2.490 ;
        RECT  3.655 0.990 3.755 1.235 ;
        RECT  3.655 1.880 3.695 2.150 ;
        RECT  3.495 0.990 3.655 2.150 ;
        RECT  3.435 1.890 3.495 2.150 ;
        RECT  3.185 0.650 3.315 0.930 ;
        RECT  3.155 0.650 3.185 2.490 ;
        RECT  3.025 0.770 3.155 2.490 ;
        RECT  2.015 0.770 3.025 0.930 ;
        RECT  2.925 1.860 3.025 2.490 ;
        RECT  2.825 0.310 2.985 0.590 ;
        RECT  2.165 1.860 2.925 2.020 ;
        RECT  2.245 1.355 2.845 1.615 ;
        RECT  1.285 0.430 2.825 0.590 ;
        RECT  1.765 1.405 2.245 1.565 ;
        RECT  2.005 1.860 2.165 2.460 ;
        RECT  1.905 2.200 2.005 2.460 ;
        RECT  1.605 0.770 1.765 1.950 ;
        RECT  1.505 0.770 1.605 0.930 ;
        RECT  1.505 1.690 1.605 1.950 ;
        RECT  1.125 0.430 1.285 2.030 ;
        RECT  0.785 0.720 1.125 0.880 ;
        RECT  0.785 1.870 1.125 2.030 ;
        RECT  0.525 0.620 0.785 0.880 ;
        RECT  0.525 1.870 0.785 2.130 ;
    END
END ADDFHX2MTH

MACRO ADDFHX4MTH
    CLASS CORE ;
    FOREIGN ADDFHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.140 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.990 1.290 22.040 1.580 ;
        RECT  21.830 0.670 21.990 2.350 ;
        RECT  21.475 0.670 21.830 0.830 ;
        RECT  21.475 2.190 21.830 2.350 ;
        RECT  21.215 0.570 21.475 0.830 ;
        RECT  21.215 2.190 21.475 2.450 ;
        END
        AntennaDiffArea 0.582 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.490 1.010 21.650 1.950 ;
        RECT  20.455 1.010 21.490 1.170 ;
        RECT  20.455 1.790 21.490 1.950 ;
        RECT  20.190 0.570 20.455 1.170 ;
        RECT  20.195 1.790 20.455 2.390 ;
        END
        AntennaDiffArea 0.573 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.370 0.880 19.580 1.170 ;
        RECT  18.905 1.010 19.370 1.170 ;
        RECT  18.645 1.010 18.905 1.330 ;
        END
        AntennaGateArea 0.4693 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.380 1.450 11.625 1.710 ;
        RECT  11.170 1.290 11.380 1.710 ;
        RECT  11.025 1.450 11.170 1.710 ;
        END
        AntennaGateArea 1.417 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.230 1.410 1.490 ;
        RECT  0.920 1.230 1.130 1.580 ;
        RECT  0.470 1.230 0.920 1.490 ;
        END
        AntennaGateArea 0.7956 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.015 -0.130 22.140 0.130 ;
        RECT  21.755 -0.130 22.015 0.490 ;
        RECT  20.965 -0.130 21.755 0.130 ;
        RECT  20.705 -0.130 20.965 0.830 ;
        RECT  19.945 -0.130 20.705 0.130 ;
        RECT  19.685 -0.130 19.945 0.670 ;
        RECT  18.895 -0.130 19.685 0.130 ;
        RECT  18.635 -0.130 18.895 0.300 ;
        RECT  13.245 -0.130 18.635 0.130 ;
        RECT  12.305 -0.130 13.245 0.250 ;
        RECT  11.485 -0.130 12.305 0.130 ;
        RECT  11.225 -0.130 11.485 0.250 ;
        RECT  1.945 -0.130 11.225 0.130 ;
        RECT  1.685 -0.130 1.945 0.250 ;
        RECT  0.895 -0.130 1.685 0.130 ;
        RECT  0.635 -0.130 0.895 0.640 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  22.015 2.740 22.140 3.000 ;
        RECT  21.755 2.530 22.015 3.000 ;
        RECT  20.965 2.740 21.755 3.000 ;
        RECT  20.705 2.230 20.965 3.000 ;
        RECT  19.845 2.740 20.705 3.000 ;
        RECT  19.245 2.620 19.845 3.000 ;
        RECT  18.325 2.740 19.245 3.000 ;
        RECT  17.385 2.620 18.325 3.000 ;
        RECT  13.475 2.740 17.385 3.000 ;
        RECT  13.215 2.570 13.475 3.000 ;
        RECT  12.425 2.740 13.215 3.000 ;
        RECT  12.165 2.235 12.425 3.000 ;
        RECT  11.405 2.740 12.165 3.000 ;
        RECT  11.145 2.235 11.405 3.000 ;
        RECT  10.385 2.740 11.145 3.000 ;
        RECT  10.125 2.235 10.385 3.000 ;
        RECT  0.895 2.740 10.125 3.000 ;
        RECT  0.635 2.235 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.295 1.350 21.305 1.510 ;
        RECT  19.475 1.690 19.635 2.440 ;
        RECT  15.535 2.280 19.475 2.440 ;
        RECT  19.175 0.440 19.440 0.700 ;
        RECT  19.135 1.350 19.295 2.100 ;
        RECT  18.365 0.540 19.175 0.700 ;
        RECT  16.555 1.940 19.135 2.100 ;
        RECT  18.365 1.600 18.915 1.760 ;
        RECT  18.260 0.540 18.365 1.760 ;
        RECT  18.205 0.310 18.260 1.760 ;
        RECT  18.095 0.310 18.205 1.315 ;
        RECT  15.885 0.310 18.095 0.470 ;
        RECT  17.585 1.155 18.095 1.315 ;
        RECT  16.905 1.600 18.005 1.760 ;
        RECT  16.905 0.650 17.835 0.810 ;
        RECT  17.085 1.105 17.585 1.365 ;
        RECT  16.745 0.650 16.905 1.760 ;
        RECT  16.645 0.650 16.745 0.810 ;
        RECT  16.395 1.840 16.555 2.100 ;
        RECT  16.235 0.680 16.395 2.100 ;
        RECT  16.135 0.680 16.235 0.930 ;
        RECT  15.445 0.770 16.135 0.930 ;
        RECT  15.945 1.820 16.045 2.080 ;
        RECT  15.785 1.255 15.945 2.080 ;
        RECT  15.625 0.310 15.885 0.575 ;
        RECT  15.105 1.255 15.785 1.415 ;
        RECT  14.695 0.310 15.625 0.470 ;
        RECT  15.435 1.900 15.535 2.440 ;
        RECT  15.285 0.650 15.445 0.930 ;
        RECT  15.275 1.630 15.435 2.560 ;
        RECT  15.055 0.650 15.285 0.810 ;
        RECT  14.765 1.630 15.275 1.790 ;
        RECT  14.415 2.400 15.275 2.560 ;
        RECT  14.945 0.990 15.105 1.415 ;
        RECT  14.695 2.010 14.955 2.220 ;
        RECT  14.695 0.990 14.945 1.150 ;
        RECT  14.605 1.330 14.765 1.790 ;
        RECT  14.535 0.310 14.695 1.150 ;
        RECT  13.875 2.010 14.695 2.170 ;
        RECT  14.185 1.330 14.605 1.490 ;
        RECT  13.845 1.670 14.425 1.830 ;
        RECT  14.155 2.355 14.415 2.560 ;
        RECT  14.025 0.500 14.185 1.490 ;
        RECT  13.405 2.010 13.875 2.270 ;
        RECT  13.685 0.310 13.845 1.830 ;
        RECT  13.585 0.310 13.685 0.590 ;
        RECT  8.635 0.430 13.585 0.590 ;
        RECT  13.345 0.770 13.505 1.580 ;
        RECT  13.195 1.895 13.405 2.270 ;
        RECT  8.975 0.770 13.345 0.930 ;
        RECT  12.935 1.895 13.195 2.055 ;
        RECT  11.975 1.110 13.155 1.270 ;
        RECT  12.675 1.895 12.935 2.380 ;
        RECT  11.975 1.895 12.675 2.055 ;
        RECT  11.915 1.110 11.975 2.055 ;
        RECT  11.815 1.110 11.915 2.375 ;
        RECT  11.765 1.110 11.815 1.270 ;
        RECT  11.655 1.895 11.815 2.375 ;
        RECT  10.895 1.895 11.655 2.055 ;
        RECT  10.845 1.110 10.945 1.270 ;
        RECT  10.845 1.895 10.895 2.495 ;
        RECT  10.685 1.110 10.845 2.495 ;
        RECT  10.635 1.895 10.685 2.495 ;
        RECT  9.875 1.895 10.635 2.055 ;
        RECT  9.315 1.110 10.005 1.270 ;
        RECT  9.775 1.895 9.875 2.495 ;
        RECT  9.615 1.450 9.775 2.495 ;
        RECT  9.525 1.450 9.615 1.710 ;
        RECT  9.155 1.110 9.315 2.560 ;
        RECT  5.165 2.400 9.155 2.560 ;
        RECT  8.815 0.770 8.975 2.220 ;
        RECT  6.485 2.060 8.815 2.220 ;
        RECT  8.475 0.430 8.635 1.880 ;
        RECT  8.305 0.430 8.475 0.645 ;
        RECT  7.245 1.720 8.475 1.880 ;
        RECT  8.205 0.385 8.305 0.645 ;
        RECT  8.045 0.385 8.205 0.925 ;
        RECT  6.995 1.380 8.175 1.540 ;
        RECT  7.255 0.765 8.045 0.925 ;
        RECT  7.535 0.310 7.795 0.585 ;
        RECT  6.715 0.310 7.535 0.470 ;
        RECT  6.995 0.650 7.255 0.925 ;
        RECT  6.735 1.380 6.995 1.880 ;
        RECT  6.715 1.380 6.735 1.600 ;
        RECT  6.555 0.310 6.715 1.600 ;
        RECT  6.455 0.310 6.555 0.690 ;
        RECT  5.975 1.440 6.555 1.600 ;
        RECT  6.225 1.835 6.485 2.220 ;
        RECT  5.665 0.310 6.455 0.470 ;
        RECT  5.505 2.060 6.225 2.220 ;
        RECT  6.075 0.695 6.175 0.955 ;
        RECT  5.915 0.695 6.075 1.245 ;
        RECT  5.815 1.440 5.975 1.880 ;
        RECT  4.615 1.085 5.915 1.245 ;
        RECT  5.685 1.720 5.815 1.880 ;
        RECT  5.405 0.310 5.665 0.905 ;
        RECT  5.345 1.880 5.505 2.220 ;
        RECT  3.815 0.310 5.405 0.470 ;
        RECT  4.705 1.880 5.345 2.040 ;
        RECT  5.005 2.230 5.165 2.560 ;
        RECT  4.145 0.650 5.155 0.810 ;
        RECT  4.145 2.330 5.005 2.490 ;
        RECT  4.565 1.880 4.705 2.150 ;
        RECT  4.565 0.990 4.615 1.245 ;
        RECT  4.405 0.990 4.565 2.150 ;
        RECT  4.355 0.990 4.405 1.150 ;
        RECT  3.985 0.650 4.145 2.490 ;
        RECT  3.845 0.770 3.985 1.030 ;
        RECT  3.255 1.860 3.985 2.020 ;
        RECT  3.045 0.770 3.845 0.930 ;
        RECT  3.655 0.310 3.815 0.590 ;
        RECT  3.065 1.355 3.690 1.615 ;
        RECT  1.885 0.430 3.655 0.590 ;
        RECT  3.095 1.860 3.255 2.300 ;
        RECT  2.990 2.040 3.095 2.300 ;
        RECT  2.485 1.405 3.065 1.565 ;
        RECT  2.780 0.770 3.045 1.030 ;
        RECT  2.345 0.810 2.485 2.145 ;
        RECT  2.325 0.810 2.345 2.495 ;
        RECT  2.225 0.810 2.325 0.970 ;
        RECT  2.085 1.885 2.325 2.495 ;
        RECT  1.685 0.430 1.885 1.950 ;
        RECT  1.405 0.430 1.685 0.590 ;
        RECT  1.405 1.790 1.685 1.950 ;
        RECT  1.145 0.400 1.405 1.000 ;
        RECT  1.145 1.790 1.405 2.390 ;
        RECT  0.385 0.840 1.145 1.000 ;
        RECT  0.385 1.790 1.145 1.950 ;
        RECT  0.125 0.400 0.385 1.000 ;
        RECT  0.125 1.790 0.385 2.390 ;
    END
END ADDFHX4MTH

MACRO ADDFHX8MTH
    CLASS CORE ;
    FOREIGN ADDFHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 27.470 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  26.885 1.495 26.960 2.195 ;
        RECT  26.880 1.495 26.885 2.390 ;
        RECT  26.835 0.655 26.880 2.390 ;
        RECT  26.625 0.405 26.835 2.390 ;
        RECT  26.575 0.405 26.625 2.055 ;
        RECT  26.510 0.655 26.575 2.055 ;
        RECT  25.875 0.655 26.510 1.005 ;
        RECT  25.865 1.705 26.510 2.055 ;
        RECT  25.615 0.405 25.875 1.005 ;
        RECT  25.605 1.705 25.865 2.460 ;
        END
        AntennaDiffArea 1.102 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  24.110 1.530 24.910 1.915 ;
        RECT  24.525 0.400 24.785 1.000 ;
        RECT  24.110 0.650 24.525 1.000 ;
        RECT  23.845 0.650 24.110 1.915 ;
        RECT  23.700 0.395 23.845 1.915 ;
        RECT  23.585 0.395 23.700 1.880 ;
        RECT  22.610 1.530 23.585 1.880 ;
        END
        AntennaDiffArea 1.308 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  20.810 1.165 22.345 1.425 ;
        RECT  20.600 0.880 20.810 1.425 ;
        RECT  20.385 1.165 20.600 1.425 ;
        END
        AntennaGateArea 0.9945 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.480 1.455 15.625 1.715 ;
        RECT  15.270 1.290 15.480 1.715 ;
        RECT  15.125 1.455 15.270 1.715 ;
        END
        AntennaGateArea 1.1531 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.230 2.265 1.490 ;
        RECT  0.510 1.230 0.720 1.580 ;
        RECT  0.405 1.230 0.510 1.490 ;
        END
        AntennaGateArea 1.5886 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  27.295 -0.130 27.470 0.130 ;
        RECT  27.135 -0.130 27.295 0.975 ;
        RECT  25.325 -0.130 27.135 0.130 ;
        RECT  25.065 -0.130 25.325 0.980 ;
        RECT  23.335 -0.130 25.065 0.130 ;
        RECT  23.075 -0.130 23.335 0.980 ;
        RECT  21.345 -0.130 23.075 0.130 ;
        RECT  21.085 -0.130 21.345 0.300 ;
        RECT  15.585 -0.130 21.085 0.130 ;
        RECT  15.325 -0.130 15.585 0.250 ;
        RECT  6.705 -0.130 15.325 0.130 ;
        RECT  6.445 -0.130 6.705 0.250 ;
        RECT  5.625 -0.130 6.445 0.130 ;
        RECT  5.365 -0.130 5.625 0.250 ;
        RECT  4.025 -0.130 5.365 0.130 ;
        RECT  3.765 -0.130 4.025 0.250 ;
        RECT  3.085 -0.130 3.765 0.130 ;
        RECT  2.825 -0.130 3.085 0.250 ;
        RECT  2.005 -0.130 2.825 0.130 ;
        RECT  1.745 -0.130 2.005 0.640 ;
        RECT  0.925 -0.130 1.745 0.130 ;
        RECT  0.665 -0.130 0.925 0.640 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.375 2.740 27.470 3.000 ;
        RECT  26.115 2.235 26.375 3.000 ;
        RECT  25.315 2.740 26.115 3.000 ;
        RECT  25.055 2.480 25.315 3.000 ;
        RECT  23.440 2.740 25.055 3.000 ;
        RECT  23.180 2.475 23.440 3.000 ;
        RECT  15.505 2.740 23.180 3.000 ;
        RECT  15.245 2.235 15.505 3.000 ;
        RECT  14.485 2.740 15.245 3.000 ;
        RECT  14.225 2.235 14.485 3.000 ;
        RECT  6.705 2.740 14.225 3.000 ;
        RECT  6.445 2.230 6.705 3.000 ;
        RECT  5.625 2.740 6.445 3.000 ;
        RECT  5.365 2.230 5.625 3.000 ;
        RECT  3.335 2.740 5.365 3.000 ;
        RECT  3.075 2.570 3.335 3.000 ;
        RECT  1.325 2.740 3.075 3.000 ;
        RECT  1.065 2.230 1.325 3.000 ;
        RECT  0.385 2.740 1.065 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  25.310 1.225 26.325 1.485 ;
        RECT  25.150 1.225 25.310 2.295 ;
        RECT  22.960 2.135 25.150 2.295 ;
        RECT  22.800 2.060 22.960 2.295 ;
        RECT  22.565 0.380 22.825 0.980 ;
        RECT  18.645 2.060 22.800 2.220 ;
        RECT  17.625 2.400 22.620 2.560 ;
        RECT  21.885 0.540 22.565 0.700 ;
        RECT  20.205 1.720 22.360 1.880 ;
        RECT  21.625 0.385 21.885 0.985 ;
        RECT  20.805 0.540 21.625 0.700 ;
        RECT  20.545 0.440 20.805 0.700 ;
        RECT  20.205 0.540 20.545 0.700 ;
        RECT  20.045 0.330 20.205 1.880 ;
        RECT  18.845 0.330 20.045 0.490 ;
        RECT  19.335 1.450 20.045 1.610 ;
        RECT  19.695 0.680 19.865 0.840 ;
        RECT  19.535 0.680 19.695 1.270 ;
        RECT  19.155 1.110 19.535 1.270 ;
        RECT  19.215 0.680 19.355 0.840 ;
        RECT  19.055 0.680 19.215 0.930 ;
        RECT  18.995 1.110 19.155 1.815 ;
        RECT  18.595 0.770 19.055 0.930 ;
        RECT  18.895 1.555 18.995 1.815 ;
        RECT  18.585 0.330 18.845 0.575 ;
        RECT  18.595 1.555 18.645 2.220 ;
        RECT  18.435 0.770 18.595 2.220 ;
        RECT  17.835 0.330 18.585 0.490 ;
        RECT  18.275 0.770 18.435 0.930 ;
        RECT  18.385 1.555 18.435 2.220 ;
        RECT  18.015 0.670 18.275 0.930 ;
        RECT  18.035 1.820 18.135 2.080 ;
        RECT  17.875 1.560 18.035 2.080 ;
        RECT  17.835 1.560 17.875 1.720 ;
        RECT  17.675 0.330 17.835 1.720 ;
        RECT  17.445 0.500 17.675 0.760 ;
        RECT  17.495 1.900 17.625 2.560 ;
        RECT  17.335 1.130 17.495 2.560 ;
        RECT  17.145 1.130 17.335 1.290 ;
        RECT  16.475 2.400 17.335 2.560 ;
        RECT  16.995 1.470 17.155 1.880 ;
        RECT  16.985 0.620 17.145 1.290 ;
        RECT  16.815 2.060 17.035 2.220 ;
        RECT  16.805 1.470 16.995 1.630 ;
        RECT  16.655 1.810 16.815 2.220 ;
        RECT  16.645 0.310 16.805 1.630 ;
        RECT  15.965 1.810 16.655 1.970 ;
        RECT  16.540 0.310 16.645 0.590 ;
        RECT  12.735 0.430 16.540 0.590 ;
        RECT  16.315 2.150 16.475 2.560 ;
        RECT  16.305 0.770 16.465 1.570 ;
        RECT  13.075 0.770 16.305 0.930 ;
        RECT  15.965 1.115 16.125 1.275 ;
        RECT  15.805 1.115 15.965 2.375 ;
        RECT  14.995 1.895 15.805 2.055 ;
        RECT  14.945 1.115 15.045 1.275 ;
        RECT  14.945 1.895 14.995 2.370 ;
        RECT  14.785 1.115 14.945 2.370 ;
        RECT  14.735 1.895 14.785 2.370 ;
        RECT  13.975 1.895 14.735 2.055 ;
        RECT  13.415 1.110 14.105 1.270 ;
        RECT  13.785 1.895 13.975 2.370 ;
        RECT  13.715 1.450 13.785 2.370 ;
        RECT  13.625 1.450 13.715 2.055 ;
        RECT  13.255 1.110 13.415 2.560 ;
        RECT  9.175 2.400 13.255 2.560 ;
        RECT  12.915 0.770 13.075 2.220 ;
        RECT  10.455 2.060 12.915 2.220 ;
        RECT  12.575 0.430 12.735 1.880 ;
        RECT  12.355 0.430 12.575 0.590 ;
        RECT  11.295 1.720 12.575 1.880 ;
        RECT  12.195 0.385 12.355 0.925 ;
        RECT  11.045 1.380 12.275 1.540 ;
        RECT  11.355 0.765 12.195 0.925 ;
        RECT  11.700 0.425 11.895 0.585 ;
        RECT  11.540 0.310 11.700 0.585 ;
        RECT  10.765 0.310 11.540 0.470 ;
        RECT  11.145 0.650 11.355 0.925 ;
        RECT  11.095 0.650 11.145 0.810 ;
        RECT  10.785 1.380 11.045 1.880 ;
        RECT  10.765 1.380 10.785 1.600 ;
        RECT  10.605 0.310 10.765 1.600 ;
        RECT  9.765 0.310 10.605 0.470 ;
        RECT  9.995 1.440 10.605 1.600 ;
        RECT  10.295 1.835 10.455 2.220 ;
        RECT  9.515 2.060 10.295 2.220 ;
        RECT  10.175 0.685 10.275 0.945 ;
        RECT  10.015 0.685 10.175 1.260 ;
        RECT  8.715 1.100 10.015 1.260 ;
        RECT  9.835 1.440 9.995 1.880 ;
        RECT  9.735 1.720 9.835 1.880 ;
        RECT  9.505 0.310 9.765 0.895 ;
        RECT  9.355 1.880 9.515 2.220 ;
        RECT  7.695 0.310 9.505 0.470 ;
        RECT  8.715 1.880 9.355 2.040 ;
        RECT  8.995 0.650 9.255 0.910 ;
        RECT  9.015 2.220 9.175 2.560 ;
        RECT  8.205 2.400 9.015 2.560 ;
        RECT  8.175 0.650 8.995 0.810 ;
        RECT  8.615 0.990 8.715 1.260 ;
        RECT  8.615 1.880 8.715 2.150 ;
        RECT  8.455 0.990 8.615 2.150 ;
        RECT  8.105 2.070 8.205 2.560 ;
        RECT  8.105 0.650 8.175 0.910 ;
        RECT  8.045 0.650 8.105 2.560 ;
        RECT  7.945 0.650 8.045 2.330 ;
        RECT  7.915 0.650 7.945 0.970 ;
        RECT  7.245 1.860 7.945 2.020 ;
        RECT  4.825 0.810 7.915 0.970 ;
        RECT  7.510 0.310 7.695 0.590 ;
        RECT  2.695 0.430 7.510 0.590 ;
        RECT  5.425 1.225 7.370 1.485 ;
        RECT  6.985 1.860 7.245 2.495 ;
        RECT  6.165 1.860 6.985 2.020 ;
        RECT  5.905 1.860 6.165 2.495 ;
        RECT  5.085 1.860 5.905 2.020 ;
        RECT  4.330 1.275 5.425 1.435 ;
        RECT  4.925 1.860 5.085 2.495 ;
        RECT  4.825 2.235 4.925 2.495 ;
        RECT  4.330 1.685 4.685 1.945 ;
        RECT  4.330 0.815 4.565 0.975 ;
        RECT  4.170 0.815 4.330 1.945 ;
        RECT  3.735 1.275 4.170 1.435 ;
        RECT  3.575 0.770 3.735 1.945 ;
        RECT  3.225 0.770 3.575 0.930 ;
        RECT  3.475 1.685 3.575 1.945 ;
        RECT  2.695 1.765 2.795 2.365 ;
        RECT  2.545 0.430 2.695 2.365 ;
        RECT  2.535 0.400 2.545 2.365 ;
        RECT  2.285 0.400 2.535 1.000 ;
        RECT  1.865 1.765 2.535 1.925 ;
        RECT  1.465 0.840 2.285 1.000 ;
        RECT  1.605 1.765 1.865 2.365 ;
        RECT  0.785 1.765 1.605 1.925 ;
        RECT  1.205 0.400 1.465 1.000 ;
        RECT  0.385 0.840 1.205 1.000 ;
        RECT  0.525 1.765 0.785 2.115 ;
        RECT  0.120 0.400 0.385 1.000 ;
    END
END ADDFHX8MTH

MACRO ADDFHXLMTH
    CLASS CORE ;
    FOREIGN ADDFHXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.220 0.730 11.380 2.050 ;
        RECT  11.170 0.730 11.220 1.170 ;
        RECT  11.090 1.790 11.220 2.050 ;
        RECT  11.095 0.730 11.170 0.990 ;
        END
        AntennaDiffArea 0.225 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.510 1.290 10.560 1.580 ;
        RECT  10.350 0.730 10.510 1.880 ;
        RECT  10.105 0.730 10.350 0.990 ;
        RECT  10.010 1.720 10.350 1.880 ;
        END
        AntennaDiffArea 0.254 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.160 0.880 9.330 1.635 ;
        RECT  9.120 0.880 9.160 1.170 ;
        END
        AntennaGateArea 0.0858 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.990 1.290 5.295 1.765 ;
        END
        AntennaGateArea 0.3458 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.210 0.485 1.470 ;
        RECT  0.100 1.090 0.360 1.665 ;
        END
        AntennaGateArea 0.1547 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.305 -0.130 11.480 0.130 ;
        RECT  10.465 -0.130 11.305 0.300 ;
        RECT  10.280 -0.130 10.465 0.130 ;
        RECT  9.440 -0.130 10.280 0.300 ;
        RECT  1.675 -0.130 9.440 0.130 ;
        RECT  0.735 -0.130 1.675 0.250 ;
        RECT  0.000 -0.130 0.735 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.180 2.740 11.480 3.000 ;
        RECT  10.580 2.560 11.180 3.000 ;
        RECT  5.495 2.740 10.580 3.000 ;
        RECT  5.235 2.285 5.495 3.000 ;
        RECT  1.500 2.740 5.235 3.000 ;
        RECT  0.900 2.390 1.500 3.000 ;
        RECT  0.000 2.740 0.900 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.900 1.350 11.035 1.610 ;
        RECT  10.740 1.330 10.900 2.220 ;
        RECT  8.190 2.060 10.740 2.220 ;
        RECT  6.605 2.400 10.395 2.560 ;
        RECT  9.760 0.685 9.855 0.945 ;
        RECT  9.755 0.685 9.760 1.880 ;
        RECT  9.595 0.540 9.755 1.880 ;
        RECT  9.245 0.540 9.595 0.700 ;
        RECT  9.500 1.720 9.595 1.880 ;
        RECT  9.085 0.310 9.245 0.700 ;
        RECT  7.685 0.310 9.085 0.470 ;
        RECT  8.750 0.735 8.875 0.895 ;
        RECT  8.590 0.735 8.750 1.880 ;
        RECT  8.400 1.720 8.590 1.880 ;
        RECT  8.190 0.735 8.305 0.895 ;
        RECT  8.030 0.735 8.190 2.220 ;
        RECT  7.830 1.750 8.030 2.010 ;
        RECT  7.525 0.310 7.685 0.945 ;
        RECT  7.455 0.785 7.525 0.945 ;
        RECT  7.295 0.785 7.455 1.935 ;
        RECT  7.175 1.775 7.295 1.935 ;
        RECT  6.775 0.310 7.250 0.470 ;
        RECT  7.015 1.775 7.175 2.155 ;
        RECT  6.955 0.685 7.115 1.595 ;
        RECT  6.915 1.895 7.015 2.155 ;
        RECT  6.605 1.435 6.955 1.595 ;
        RECT  6.615 0.310 6.775 1.255 ;
        RECT  3.885 0.310 6.615 0.470 ;
        RECT  6.185 1.095 6.615 1.255 ;
        RECT  6.445 1.435 6.605 2.560 ;
        RECT  6.345 2.165 6.445 2.425 ;
        RECT  6.275 0.650 6.435 0.915 ;
        RECT  5.695 0.755 6.275 0.915 ;
        RECT  6.025 1.095 6.185 1.975 ;
        RECT  5.835 2.235 6.010 2.495 ;
        RECT  5.695 1.945 5.835 2.495 ;
        RECT  5.675 0.755 5.695 2.495 ;
        RECT  5.535 0.755 5.675 2.105 ;
        RECT  4.985 1.945 5.535 2.105 ;
        RECT  5.035 0.850 5.325 1.110 ;
        RECT  4.875 0.650 5.035 1.110 ;
        RECT  4.765 1.945 4.985 2.485 ;
        RECT  4.255 0.650 4.875 0.810 ;
        RECT  4.725 1.855 4.765 2.485 ;
        RECT  4.605 1.855 4.725 2.115 ;
        RECT  4.595 0.990 4.695 1.150 ;
        RECT  4.435 0.990 4.595 1.385 ;
        RECT  4.425 1.225 4.435 1.385 ;
        RECT  4.265 1.225 4.425 2.560 ;
        RECT  2.225 2.400 4.265 2.560 ;
        RECT  4.095 0.650 4.255 1.045 ;
        RECT  4.085 0.885 4.095 1.045 ;
        RECT  3.925 0.885 4.085 2.220 ;
        RECT  2.735 2.060 3.925 2.220 ;
        RECT  3.745 0.310 3.885 0.705 ;
        RECT  3.725 0.310 3.745 1.880 ;
        RECT  3.585 0.545 3.725 1.880 ;
        RECT  3.485 1.720 3.585 1.880 ;
        RECT  3.235 0.430 3.325 1.470 ;
        RECT  3.165 0.430 3.235 1.880 ;
        RECT  0.890 0.430 3.165 0.590 ;
        RECT  3.075 1.310 3.165 1.880 ;
        RECT  2.975 1.720 3.075 1.880 ;
        RECT  2.735 0.775 2.785 0.935 ;
        RECT  2.575 0.775 2.735 2.220 ;
        RECT  2.525 0.775 2.575 0.935 ;
        RECT  2.465 1.800 2.575 2.060 ;
        RECT  2.225 0.770 2.275 0.930 ;
        RECT  2.065 0.770 2.225 2.560 ;
        RECT  2.015 0.770 2.065 0.930 ;
        RECT  1.955 1.800 2.065 2.060 ;
        RECT  1.580 1.285 1.840 1.545 ;
        RECT  1.365 1.335 1.580 1.495 ;
        RECT  1.205 0.770 1.365 1.905 ;
        RECT  1.105 0.770 1.205 0.930 ;
        RECT  1.095 1.645 1.205 1.905 ;
        RECT  0.730 0.430 0.890 2.005 ;
        RECT  0.125 0.745 0.730 0.905 ;
        RECT  0.385 1.845 0.730 2.005 ;
        RECT  0.125 1.845 0.385 2.105 ;
    END
END ADDFHXLMTH

MACRO ADDFX1MTH
    CLASS CORE ;
    FOREIGN ADDFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.485 1.700 10.560 1.990 ;
        RECT  10.325 0.685 10.485 1.990 ;
        END
        AntennaDiffArea 0.333 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.440 1.720 9.495 1.880 ;
        RECT  9.230 0.685 9.440 1.880 ;
        RECT  9.180 0.685 9.230 1.170 ;
        RECT  9.120 0.880 9.180 1.170 ;
        END
        AntennaDiffArea 0.333 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.350 1.110 7.465 1.270 ;
        RECT  7.350 1.900 7.400 2.060 ;
        RECT  7.190 1.110 7.350 2.060 ;
        RECT  7.070 1.285 7.190 1.580 ;
        RECT  7.140 1.900 7.190 2.060 ;
        END
        AntennaGateArea 0.1742 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.265 0.430 1.525 ;
        RECT  0.100 1.265 0.310 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.110 3.730 1.375 ;
        RECT  3.380 1.110 3.590 1.580 ;
        END
        AntennaGateArea 0.208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.980 -0.130 10.660 0.130 ;
        RECT  9.720 -0.130 9.980 0.675 ;
        RECT  9.090 -0.130 9.720 0.335 ;
        RECT  8.215 -0.130 9.090 0.130 ;
        RECT  7.275 -0.130 8.215 0.250 ;
        RECT  3.535 -0.130 7.275 0.130 ;
        RECT  3.245 -0.130 3.535 0.250 ;
        RECT  0.895 -0.130 3.245 0.130 ;
        RECT  0.635 -0.130 0.895 0.625 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 2.740 10.660 3.000 ;
        RECT  9.805 2.555 10.405 3.000 ;
        RECT  7.320 2.740 9.805 3.000 ;
        RECT  7.060 2.620 7.320 3.000 ;
        RECT  3.615 2.740 7.060 3.000 ;
        RECT  3.355 2.620 3.615 3.000 ;
        RECT  0.925 2.740 3.355 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.985 1.175 10.145 1.435 ;
        RECT  9.875 1.275 9.985 1.435 ;
        RECT  9.715 1.275 9.875 2.220 ;
        RECT  8.355 2.060 9.715 2.220 ;
        RECT  7.665 2.400 9.595 2.560 ;
        RECT  8.880 1.705 8.985 1.865 ;
        RECT  8.720 0.430 8.880 1.865 ;
        RECT  6.990 0.430 8.720 0.590 ;
        RECT  8.355 0.770 8.420 0.930 ;
        RECT  8.195 0.770 8.355 2.220 ;
        RECT  8.160 0.770 8.195 0.930 ;
        RECT  7.765 0.770 7.925 2.060 ;
        RECT  6.610 0.770 7.765 0.930 ;
        RECT  7.685 1.800 7.765 2.060 ;
        RECT  7.505 2.280 7.665 2.560 ;
        RECT  6.885 2.280 7.505 2.440 ;
        RECT  6.830 0.310 6.990 0.590 ;
        RECT  6.725 2.280 6.885 2.545 ;
        RECT  6.710 1.110 6.870 1.850 ;
        RECT  4.775 0.310 6.830 0.470 ;
        RECT  6.105 2.385 6.725 2.545 ;
        RECT  6.610 1.110 6.710 1.270 ;
        RECT  6.545 1.690 6.710 1.850 ;
        RECT  6.445 0.670 6.610 0.930 ;
        RECT  6.385 1.690 6.545 2.205 ;
        RECT  5.305 0.670 6.445 0.830 ;
        RECT  6.285 2.045 6.385 2.205 ;
        RECT  6.105 1.110 6.270 1.270 ;
        RECT  5.945 1.110 6.105 2.545 ;
        RECT  5.585 2.290 5.945 2.545 ;
        RECT  5.605 1.110 5.765 2.100 ;
        RECT  5.485 1.110 5.605 1.270 ;
        RECT  5.335 1.940 5.605 2.100 ;
        RECT  5.305 1.500 5.425 1.760 ;
        RECT  5.175 1.940 5.335 2.440 ;
        RECT  5.145 0.670 5.305 1.760 ;
        RECT  5.075 2.225 5.175 2.440 ;
        RECT  4.740 1.600 5.145 1.760 ;
        RECT  4.425 2.280 5.075 2.440 ;
        RECT  4.315 1.260 4.965 1.420 ;
        RECT  4.615 0.310 4.775 0.875 ;
        RECT  4.580 1.600 4.740 2.100 ;
        RECT  3.875 0.310 4.615 0.470 ;
        RECT  2.605 1.940 4.580 2.100 ;
        RECT  4.165 2.280 4.425 2.545 ;
        RECT  4.155 0.665 4.315 1.760 ;
        RECT  2.620 2.280 4.165 2.440 ;
        RECT  4.055 0.665 4.155 0.930 ;
        RECT  3.935 1.600 4.155 1.760 ;
        RECT  2.805 0.770 4.055 0.930 ;
        RECT  3.715 0.310 3.875 0.590 ;
        RECT  3.055 0.430 3.715 0.590 ;
        RECT  2.895 0.325 3.055 0.590 ;
        RECT  2.945 1.600 3.045 1.760 ;
        RECT  2.805 1.155 2.945 1.760 ;
        RECT  1.765 0.325 2.895 0.485 ;
        RECT  2.785 0.770 2.805 1.760 ;
        RECT  2.715 0.770 2.785 1.315 ;
        RECT  2.645 0.665 2.715 1.315 ;
        RECT  2.455 0.665 2.645 0.930 ;
        RECT  2.460 2.280 2.620 2.545 ;
        RECT  2.445 1.585 2.605 2.100 ;
        RECT  1.260 2.385 2.460 2.545 ;
        RECT  2.380 1.585 2.445 1.745 ;
        RECT  2.220 1.150 2.380 1.745 ;
        RECT  1.600 2.045 2.265 2.205 ;
        RECT  2.205 1.150 2.220 1.310 ;
        RECT  2.045 0.665 2.205 1.310 ;
        RECT  1.945 0.665 2.045 0.825 ;
        RECT  1.765 1.600 2.040 1.760 ;
        RECT  1.605 0.325 1.765 1.760 ;
        RECT  1.440 1.940 1.600 2.205 ;
        RECT  1.355 1.940 1.440 2.100 ;
        RECT  1.195 0.615 1.355 2.100 ;
        RECT  1.100 2.280 1.260 2.545 ;
        RECT  0.985 2.280 1.100 2.440 ;
        RECT  0.825 0.865 0.985 2.440 ;
        RECT  0.335 0.865 0.825 1.025 ;
        RECT  0.335 2.280 0.825 2.440 ;
        RECT  0.175 0.425 0.335 1.025 ;
        RECT  0.175 2.170 0.335 2.440 ;
    END
END ADDFX1MTH

MACRO ADDFX2MTH
    CLASS CORE ;
    FOREIGN ADDFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.300 0.345 10.560 2.285 ;
        END
        AntennaDiffArea 0.527 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.185 0.345 9.445 1.875 ;
        RECT  9.120 0.880 9.185 1.170 ;
        END
        AntennaDiffArea 0.521 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.300 1.110 7.415 1.270 ;
        RECT  7.300 1.900 7.350 2.060 ;
        RECT  7.140 1.110 7.300 2.060 ;
        RECT  7.070 1.285 7.140 1.580 ;
        RECT  7.090 1.900 7.140 2.060 ;
        END
        AntennaGateArea 0.1742 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.265 0.450 1.525 ;
        RECT  0.100 1.265 0.310 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.110 3.680 1.375 ;
        RECT  3.380 1.110 3.590 1.580 ;
        END
        AntennaGateArea 0.208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.995 -0.130 10.660 0.130 ;
        RECT  9.735 -0.130 9.995 0.955 ;
        RECT  8.760 -0.130 9.735 0.130 ;
        RECT  8.500 -0.130 8.760 0.250 ;
        RECT  8.165 -0.130 8.500 0.130 ;
        RECT  7.225 -0.130 8.165 0.250 ;
        RECT  3.485 -0.130 7.225 0.130 ;
        RECT  3.195 -0.130 3.485 0.250 ;
        RECT  0.905 -0.130 3.195 0.130 ;
        RECT  0.645 -0.130 0.905 0.625 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.990 2.740 10.660 3.000 ;
        RECT  9.730 2.415 9.990 3.000 ;
        RECT  7.270 2.740 9.730 3.000 ;
        RECT  7.010 2.620 7.270 3.000 ;
        RECT  3.565 2.740 7.010 3.000 ;
        RECT  3.305 2.620 3.565 3.000 ;
        RECT  0.925 2.740 3.305 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.920 1.175 10.080 2.220 ;
        RECT  8.305 2.060 9.920 2.220 ;
        RECT  7.615 2.400 9.125 2.560 ;
        RECT  8.890 1.705 8.935 1.865 ;
        RECT  8.730 0.430 8.890 1.865 ;
        RECT  6.940 0.430 8.730 0.590 ;
        RECT  8.675 1.705 8.730 1.865 ;
        RECT  8.305 0.770 8.430 0.930 ;
        RECT  8.145 0.770 8.305 2.220 ;
        RECT  7.855 0.770 7.920 0.930 ;
        RECT  7.695 0.770 7.855 2.060 ;
        RECT  6.560 0.770 7.695 0.930 ;
        RECT  7.635 1.800 7.695 2.060 ;
        RECT  7.455 2.240 7.615 2.560 ;
        RECT  6.835 2.240 7.455 2.400 ;
        RECT  6.780 0.310 6.940 0.590 ;
        RECT  6.675 2.240 6.835 2.545 ;
        RECT  6.660 1.110 6.820 1.850 ;
        RECT  4.725 0.310 6.780 0.470 ;
        RECT  6.055 2.385 6.675 2.545 ;
        RECT  6.560 1.110 6.660 1.270 ;
        RECT  6.495 1.690 6.660 1.850 ;
        RECT  6.395 0.670 6.560 0.930 ;
        RECT  6.335 1.690 6.495 2.205 ;
        RECT  5.255 0.670 6.395 0.830 ;
        RECT  6.235 2.045 6.335 2.205 ;
        RECT  6.055 1.110 6.220 1.270 ;
        RECT  5.895 1.110 6.055 2.545 ;
        RECT  5.535 2.290 5.895 2.545 ;
        RECT  5.555 1.110 5.715 2.100 ;
        RECT  5.435 1.110 5.555 1.270 ;
        RECT  5.285 1.940 5.555 2.100 ;
        RECT  5.255 1.500 5.375 1.760 ;
        RECT  5.125 1.940 5.285 2.440 ;
        RECT  5.095 0.670 5.255 1.760 ;
        RECT  5.025 2.225 5.125 2.440 ;
        RECT  4.690 1.600 5.095 1.760 ;
        RECT  4.375 2.280 5.025 2.440 ;
        RECT  4.265 1.260 4.915 1.420 ;
        RECT  4.565 0.310 4.725 0.875 ;
        RECT  4.530 1.600 4.690 2.100 ;
        RECT  3.825 0.310 4.565 0.470 ;
        RECT  2.555 1.940 4.530 2.100 ;
        RECT  4.115 2.280 4.375 2.545 ;
        RECT  4.105 0.665 4.265 1.760 ;
        RECT  2.570 2.280 4.115 2.440 ;
        RECT  4.005 0.665 4.105 0.930 ;
        RECT  3.885 1.600 4.105 1.760 ;
        RECT  2.755 0.770 4.005 0.930 ;
        RECT  3.665 0.310 3.825 0.590 ;
        RECT  3.005 0.430 3.665 0.590 ;
        RECT  2.845 0.325 3.005 0.590 ;
        RECT  2.895 1.600 2.995 1.760 ;
        RECT  2.755 1.155 2.895 1.760 ;
        RECT  1.715 0.325 2.845 0.485 ;
        RECT  2.735 0.770 2.755 1.760 ;
        RECT  2.665 0.770 2.735 1.315 ;
        RECT  2.595 0.665 2.665 1.315 ;
        RECT  2.405 0.665 2.595 0.930 ;
        RECT  2.410 2.280 2.570 2.545 ;
        RECT  2.395 1.585 2.555 2.100 ;
        RECT  1.310 2.385 2.410 2.545 ;
        RECT  2.330 1.585 2.395 1.745 ;
        RECT  2.170 1.150 2.330 1.745 ;
        RECT  1.650 2.045 2.215 2.205 ;
        RECT  2.155 1.150 2.170 1.310 ;
        RECT  1.995 0.665 2.155 1.310 ;
        RECT  1.895 0.665 1.995 0.825 ;
        RECT  1.830 1.575 1.990 1.835 ;
        RECT  1.715 1.575 1.830 1.735 ;
        RECT  1.555 0.325 1.715 1.735 ;
        RECT  1.490 1.940 1.650 2.205 ;
        RECT  1.375 1.940 1.490 2.100 ;
        RECT  1.215 0.615 1.375 2.100 ;
        RECT  1.150 2.280 1.310 2.545 ;
        RECT  1.005 2.280 1.150 2.440 ;
        RECT  0.845 0.865 1.005 2.440 ;
        RECT  0.335 0.865 0.845 1.025 ;
        RECT  0.335 2.280 0.845 2.440 ;
        RECT  0.175 0.425 0.335 1.025 ;
        RECT  0.175 2.170 0.335 2.440 ;
    END
END ADDFX2MTH

MACRO ADDFX4MTH
    CLASS CORE ;
    FOREIGN ADDFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.855 1.290 10.970 1.580 ;
        RECT  10.635 0.355 10.855 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.765 0.355 9.825 0.955 ;
        RECT  9.505 0.355 9.765 1.895 ;
        END
        AntennaDiffArea 0.596 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 1.110 7.305 2.060 ;
        END
        AntennaGateArea 0.1742 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.265 0.430 1.575 ;
        RECT  0.100 1.265 0.310 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.110 3.725 1.375 ;
        RECT  3.380 1.110 3.590 1.580 ;
        END
        AntennaGateArea 0.208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 -0.130 11.480 0.130 ;
        RECT  11.095 -0.130 11.355 1.025 ;
        RECT  10.335 -0.130 11.095 0.130 ;
        RECT  10.075 -0.130 10.335 0.955 ;
        RECT  9.315 -0.130 10.075 0.130 ;
        RECT  9.055 -0.130 9.315 0.955 ;
        RECT  8.705 -0.130 9.055 0.130 ;
        RECT  8.105 -0.130 8.705 0.250 ;
        RECT  7.740 -0.130 8.105 0.130 ;
        RECT  7.140 -0.130 7.740 0.250 ;
        RECT  3.505 -0.130 7.140 0.130 ;
        RECT  3.245 -0.130 3.505 0.250 ;
        RECT  0.915 -0.130 3.245 0.130 ;
        RECT  0.655 -0.130 0.915 0.720 ;
        RECT  0.000 -0.130 0.655 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 2.740 11.480 3.000 ;
        RECT  11.095 1.915 11.355 3.000 ;
        RECT  10.305 2.740 11.095 3.000 ;
        RECT  10.045 2.430 10.305 3.000 ;
        RECT  7.165 2.740 10.045 3.000 ;
        RECT  6.905 2.620 7.165 3.000 ;
        RECT  3.525 2.740 6.905 3.000 ;
        RECT  3.265 2.620 3.525 3.000 ;
        RECT  0.925 2.740 3.265 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.330 1.175 10.425 1.435 ;
        RECT  10.170 1.175 10.330 2.250 ;
        RECT  9.315 2.090 10.170 2.250 ;
        RECT  9.155 2.060 9.315 2.250 ;
        RECT  8.205 2.060 9.155 2.220 ;
        RECT  7.715 2.400 8.995 2.560 ;
        RECT  8.755 1.720 8.795 1.880 ;
        RECT  8.595 0.430 8.755 1.880 ;
        RECT  6.960 0.430 8.595 0.590 ;
        RECT  8.535 1.720 8.595 1.880 ;
        RECT  8.205 0.770 8.295 0.930 ;
        RECT  8.045 0.770 8.205 2.220 ;
        RECT  7.965 0.770 8.045 0.930 ;
        RECT  7.685 0.770 7.785 0.930 ;
        RECT  7.685 1.940 7.745 2.100 ;
        RECT  7.555 2.280 7.715 2.560 ;
        RECT  7.525 0.770 7.685 2.100 ;
        RECT  6.735 2.280 7.555 2.440 ;
        RECT  6.455 0.770 7.525 0.930 ;
        RECT  7.485 1.940 7.525 2.100 ;
        RECT  6.800 0.310 6.960 0.590 ;
        RECT  4.815 0.310 6.800 0.470 ;
        RECT  6.615 1.110 6.775 1.850 ;
        RECT  6.575 2.280 6.735 2.560 ;
        RECT  6.505 1.110 6.615 1.270 ;
        RECT  6.415 1.690 6.615 1.850 ;
        RECT  5.975 2.400 6.575 2.560 ;
        RECT  6.290 0.715 6.455 0.930 ;
        RECT  6.255 1.690 6.415 2.190 ;
        RECT  5.275 0.715 6.290 0.875 ;
        RECT  6.155 2.030 6.255 2.190 ;
        RECT  5.975 1.110 6.175 1.270 ;
        RECT  5.815 1.110 5.975 2.560 ;
        RECT  5.455 2.290 5.815 2.560 ;
        RECT  5.475 1.060 5.635 2.110 ;
        RECT  5.455 1.060 5.475 1.320 ;
        RECT  5.205 1.950 5.475 2.110 ;
        RECT  5.275 1.510 5.295 1.770 ;
        RECT  5.115 0.715 5.275 1.770 ;
        RECT  5.045 1.950 5.205 2.440 ;
        RECT  4.610 1.610 5.115 1.770 ;
        RECT  4.370 2.280 5.045 2.440 ;
        RECT  4.775 1.040 4.935 1.420 ;
        RECT  4.555 0.310 4.815 0.825 ;
        RECT  4.270 1.260 4.775 1.420 ;
        RECT  4.450 1.610 4.610 2.100 ;
        RECT  3.845 0.310 4.555 0.470 ;
        RECT  2.605 1.940 4.450 2.100 ;
        RECT  4.110 2.280 4.370 2.545 ;
        RECT  4.110 0.665 4.270 1.760 ;
        RECT  4.010 0.665 4.110 0.930 ;
        RECT  3.805 1.600 4.110 1.760 ;
        RECT  2.620 2.280 4.110 2.440 ;
        RECT  2.775 0.770 4.010 0.930 ;
        RECT  3.685 0.310 3.845 0.590 ;
        RECT  3.010 0.430 3.685 0.590 ;
        RECT  2.945 1.600 3.045 1.760 ;
        RECT  2.850 0.310 3.010 0.590 ;
        RECT  2.785 1.250 2.945 1.760 ;
        RECT  1.735 0.310 2.850 0.470 ;
        RECT  2.775 1.250 2.785 1.410 ;
        RECT  2.685 0.770 2.775 1.410 ;
        RECT  2.615 0.665 2.685 1.410 ;
        RECT  2.460 2.280 2.620 2.545 ;
        RECT  2.425 0.665 2.615 0.930 ;
        RECT  2.445 1.610 2.605 2.100 ;
        RECT  1.260 2.385 2.460 2.545 ;
        RECT  2.435 1.610 2.445 1.770 ;
        RECT  2.275 1.150 2.435 1.770 ;
        RECT  2.175 1.150 2.275 1.310 ;
        RECT  1.640 2.045 2.265 2.205 ;
        RECT  2.015 0.665 2.175 1.310 ;
        RECT  1.890 1.575 2.050 1.835 ;
        RECT  1.915 0.665 2.015 0.825 ;
        RECT  1.735 1.575 1.890 1.735 ;
        RECT  1.575 0.310 1.735 1.735 ;
        RECT  1.480 1.940 1.640 2.205 ;
        RECT  1.395 1.940 1.480 2.100 ;
        RECT  1.235 0.615 1.395 2.100 ;
        RECT  1.100 2.280 1.260 2.545 ;
        RECT  1.025 2.280 1.100 2.440 ;
        RECT  0.865 0.920 1.025 2.440 ;
        RECT  0.385 0.920 0.865 1.080 ;
        RECT  0.385 2.280 0.865 2.440 ;
        RECT  0.125 0.425 0.385 1.080 ;
        RECT  0.125 2.180 0.385 2.440 ;
    END
END ADDFX4MTH

MACRO ADDFX8MTH
    CLASS CORE ;
    FOREIGN ADDFX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.635 0.355 12.895 2.285 ;
        RECT  11.875 1.085 12.635 1.785 ;
        RECT  11.615 0.355 11.875 2.285 ;
        END
        AntennaDiffArea 1.2 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 0.355 10.795 1.895 ;
        RECT  9.775 1.085 10.535 1.785 ;
        RECT  9.515 0.355 9.775 1.895 ;
        RECT  9.395 1.735 9.515 1.895 ;
        END
        AntennaDiffArea 1.192 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.255 1.110 7.295 1.580 ;
        RECT  6.995 1.110 7.255 2.060 ;
        END
        AntennaGateArea 0.1742 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.265 0.430 1.575 ;
        RECT  0.100 1.265 0.310 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.110 3.695 1.375 ;
        RECT  3.380 1.110 3.590 1.580 ;
        END
        AntennaGateArea 0.208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 -0.130 13.530 0.130 ;
        RECT  13.145 -0.130 13.405 1.025 ;
        RECT  12.385 -0.130 13.145 0.130 ;
        RECT  12.125 -0.130 12.385 0.820 ;
        RECT  11.315 -0.130 12.125 0.130 ;
        RECT  11.055 -0.130 11.315 0.955 ;
        RECT  10.285 -0.130 11.055 0.130 ;
        RECT  10.025 -0.130 10.285 0.905 ;
        RECT  9.265 -0.130 10.025 0.130 ;
        RECT  9.005 -0.130 9.265 0.955 ;
        RECT  8.675 -0.130 9.005 0.130 ;
        RECT  8.075 -0.130 8.675 0.250 ;
        RECT  7.710 -0.130 8.075 0.130 ;
        RECT  7.110 -0.130 7.710 0.250 ;
        RECT  3.475 -0.130 7.110 0.130 ;
        RECT  3.215 -0.130 3.475 0.250 ;
        RECT  0.910 -0.130 3.215 0.130 ;
        RECT  0.640 -0.130 0.910 0.720 ;
        RECT  0.000 -0.130 0.640 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.915 13.405 3.000 ;
        RECT  12.385 2.740 13.145 3.000 ;
        RECT  12.125 1.965 12.385 3.000 ;
        RECT  11.335 2.740 12.125 3.000 ;
        RECT  11.075 2.445 11.335 3.000 ;
        RECT  10.255 2.740 11.075 3.000 ;
        RECT  9.995 2.445 10.255 3.000 ;
        RECT  7.115 2.740 9.995 3.000 ;
        RECT  6.855 2.620 7.115 3.000 ;
        RECT  3.515 2.740 6.855 3.000 ;
        RECT  3.255 2.620 3.515 3.000 ;
        RECT  0.925 2.740 3.255 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.245 1.160 11.405 2.265 ;
        RECT  9.265 2.105 11.245 2.265 ;
        RECT  9.105 2.060 9.265 2.265 ;
        RECT  8.155 2.060 9.105 2.220 ;
        RECT  7.665 2.400 8.945 2.560 ;
        RECT  8.705 1.720 8.745 1.880 ;
        RECT  8.545 0.430 8.705 1.880 ;
        RECT  6.930 0.430 8.545 0.590 ;
        RECT  8.485 1.720 8.545 1.880 ;
        RECT  8.155 0.770 8.305 0.930 ;
        RECT  7.995 0.770 8.155 2.220 ;
        RECT  7.915 0.770 7.995 0.930 ;
        RECT  7.655 0.770 7.735 0.930 ;
        RECT  7.655 1.940 7.695 2.100 ;
        RECT  7.505 2.280 7.665 2.560 ;
        RECT  7.495 0.770 7.655 2.100 ;
        RECT  6.685 2.280 7.505 2.440 ;
        RECT  6.425 0.770 7.495 0.930 ;
        RECT  7.435 1.940 7.495 2.100 ;
        RECT  6.770 0.310 6.930 0.590 ;
        RECT  5.915 0.310 6.770 0.470 ;
        RECT  6.585 1.110 6.745 1.850 ;
        RECT  6.525 2.280 6.685 2.560 ;
        RECT  6.475 1.110 6.585 1.270 ;
        RECT  6.365 1.690 6.585 1.850 ;
        RECT  5.925 2.400 6.525 2.560 ;
        RECT  6.260 0.715 6.425 0.930 ;
        RECT  6.205 1.690 6.365 2.190 ;
        RECT  5.225 0.715 6.260 0.875 ;
        RECT  6.105 2.030 6.205 2.190 ;
        RECT  5.925 1.110 6.125 1.270 ;
        RECT  5.765 1.110 5.925 2.560 ;
        RECT  5.655 0.310 5.915 0.490 ;
        RECT  5.415 2.290 5.765 2.560 ;
        RECT  4.775 0.310 5.655 0.470 ;
        RECT  5.405 1.060 5.565 2.110 ;
        RECT  5.155 1.950 5.405 2.110 ;
        RECT  5.065 0.715 5.225 1.770 ;
        RECT  4.995 1.950 5.155 2.440 ;
        RECT  4.545 1.610 5.065 1.770 ;
        RECT  4.330 2.280 4.995 2.440 ;
        RECT  4.680 1.040 4.840 1.420 ;
        RECT  4.515 0.310 4.775 0.825 ;
        RECT  4.200 1.260 4.680 1.420 ;
        RECT  4.385 1.610 4.545 2.100 ;
        RECT  3.815 0.310 4.515 0.470 ;
        RECT  2.575 1.940 4.385 2.100 ;
        RECT  4.070 2.280 4.330 2.545 ;
        RECT  4.200 0.665 4.240 0.825 ;
        RECT  4.040 0.665 4.200 1.760 ;
        RECT  2.590 2.280 4.070 2.440 ;
        RECT  3.980 0.665 4.040 0.930 ;
        RECT  3.795 1.600 4.040 1.760 ;
        RECT  2.745 0.770 3.980 0.930 ;
        RECT  3.655 0.310 3.815 0.590 ;
        RECT  2.980 0.430 3.655 0.590 ;
        RECT  2.915 1.600 3.015 1.760 ;
        RECT  2.820 0.310 2.980 0.590 ;
        RECT  2.755 1.250 2.915 1.760 ;
        RECT  1.705 0.310 2.820 0.470 ;
        RECT  2.745 1.250 2.755 1.410 ;
        RECT  2.655 0.770 2.745 1.410 ;
        RECT  2.585 0.665 2.655 1.410 ;
        RECT  2.430 2.280 2.590 2.545 ;
        RECT  2.395 0.665 2.585 0.930 ;
        RECT  2.415 1.610 2.575 2.100 ;
        RECT  1.260 2.385 2.430 2.545 ;
        RECT  2.405 1.610 2.415 1.770 ;
        RECT  2.245 1.150 2.405 1.770 ;
        RECT  2.145 1.150 2.245 1.310 ;
        RECT  1.610 2.045 2.235 2.205 ;
        RECT  1.985 0.665 2.145 1.310 ;
        RECT  1.860 1.575 2.020 1.835 ;
        RECT  1.885 0.665 1.985 0.825 ;
        RECT  1.705 1.575 1.860 1.735 ;
        RECT  1.545 0.310 1.705 1.735 ;
        RECT  1.450 1.940 1.610 2.205 ;
        RECT  1.365 1.940 1.450 2.100 ;
        RECT  1.205 0.615 1.365 2.100 ;
        RECT  1.100 2.280 1.260 2.545 ;
        RECT  0.995 2.280 1.100 2.440 ;
        RECT  0.835 0.920 0.995 2.440 ;
        RECT  0.385 0.920 0.835 1.080 ;
        RECT  0.385 2.280 0.835 2.440 ;
        RECT  0.125 0.425 0.385 1.080 ;
        RECT  0.125 2.180 0.385 2.440 ;
    END
END ADDFX8MTH

MACRO ADDFXLMTH
    CLASS CORE ;
    FOREIGN ADDFXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.485 1.700 10.560 1.990 ;
        RECT  10.325 0.685 10.485 1.990 ;
        END
        AntennaDiffArea 0.225 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.440 1.720 9.495 1.880 ;
        RECT  9.230 0.685 9.440 1.880 ;
        RECT  9.180 0.685 9.230 1.170 ;
        RECT  9.120 0.880 9.180 1.170 ;
        END
        AntennaDiffArea 0.229 ;
    END CO
    PIN CI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.350 1.110 7.465 1.270 ;
        RECT  7.350 1.900 7.400 2.060 ;
        RECT  7.190 1.110 7.350 2.060 ;
        RECT  7.070 1.285 7.190 1.580 ;
        RECT  7.140 1.900 7.190 2.060 ;
        END
        AntennaGateArea 0.1742 ;
    END CI
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.265 0.430 1.525 ;
        RECT  0.100 1.265 0.310 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.110 3.730 1.375 ;
        RECT  3.380 1.110 3.590 1.580 ;
        END
        AntennaGateArea 0.208 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.965 -0.130 10.660 0.130 ;
        RECT  9.705 -0.130 9.965 0.360 ;
        RECT  7.535 -0.130 9.705 0.130 ;
        RECT  7.275 -0.130 7.535 0.250 ;
        RECT  3.535 -0.130 7.275 0.130 ;
        RECT  3.245 -0.130 3.535 0.250 ;
        RECT  0.895 -0.130 3.245 0.130 ;
        RECT  0.635 -0.130 0.895 0.625 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.035 2.740 10.660 3.000 ;
        RECT  9.775 2.415 10.035 3.000 ;
        RECT  7.320 2.740 9.775 3.000 ;
        RECT  7.060 2.620 7.320 3.000 ;
        RECT  3.615 2.740 7.060 3.000 ;
        RECT  3.355 2.620 3.615 3.000 ;
        RECT  0.925 2.740 3.355 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.985 1.175 10.145 1.435 ;
        RECT  9.875 1.275 9.985 1.435 ;
        RECT  9.715 1.275 9.875 2.220 ;
        RECT  8.355 2.060 9.715 2.220 ;
        RECT  7.665 2.400 9.490 2.560 ;
        RECT  8.880 1.705 8.985 1.865 ;
        RECT  8.720 0.430 8.880 1.865 ;
        RECT  6.990 0.430 8.720 0.590 ;
        RECT  8.355 0.770 8.435 0.930 ;
        RECT  8.195 0.770 8.355 2.220 ;
        RECT  8.115 0.770 8.195 0.930 ;
        RECT  7.750 0.770 7.910 2.060 ;
        RECT  6.610 0.770 7.750 0.930 ;
        RECT  7.635 1.800 7.750 2.060 ;
        RECT  7.505 2.280 7.665 2.560 ;
        RECT  6.885 2.280 7.505 2.440 ;
        RECT  6.830 0.310 6.990 0.590 ;
        RECT  6.725 2.280 6.885 2.545 ;
        RECT  6.710 1.110 6.870 1.850 ;
        RECT  4.775 0.310 6.830 0.470 ;
        RECT  6.105 2.385 6.725 2.545 ;
        RECT  6.610 1.110 6.710 1.270 ;
        RECT  6.545 1.690 6.710 1.850 ;
        RECT  6.445 0.670 6.610 0.930 ;
        RECT  6.385 1.690 6.545 2.205 ;
        RECT  5.305 0.670 6.445 0.830 ;
        RECT  6.285 2.045 6.385 2.205 ;
        RECT  6.105 1.110 6.270 1.270 ;
        RECT  5.945 1.110 6.105 2.545 ;
        RECT  5.585 2.290 5.945 2.545 ;
        RECT  5.605 1.110 5.765 2.100 ;
        RECT  5.485 1.110 5.605 1.270 ;
        RECT  5.335 1.940 5.605 2.100 ;
        RECT  5.305 1.500 5.425 1.760 ;
        RECT  5.175 1.940 5.335 2.440 ;
        RECT  5.145 0.670 5.305 1.760 ;
        RECT  5.075 2.225 5.175 2.440 ;
        RECT  4.740 1.600 5.145 1.760 ;
        RECT  4.425 2.280 5.075 2.440 ;
        RECT  4.315 1.260 4.965 1.420 ;
        RECT  4.615 0.310 4.775 0.875 ;
        RECT  4.580 1.600 4.740 2.100 ;
        RECT  3.875 0.310 4.615 0.470 ;
        RECT  2.605 1.940 4.580 2.100 ;
        RECT  4.165 2.280 4.425 2.545 ;
        RECT  4.155 0.665 4.315 1.760 ;
        RECT  2.620 2.280 4.165 2.440 ;
        RECT  4.055 0.665 4.155 0.930 ;
        RECT  3.935 1.600 4.155 1.760 ;
        RECT  2.805 0.770 4.055 0.930 ;
        RECT  3.715 0.310 3.875 0.590 ;
        RECT  3.055 0.430 3.715 0.590 ;
        RECT  2.895 0.325 3.055 0.590 ;
        RECT  2.945 1.600 3.045 1.760 ;
        RECT  2.805 1.155 2.945 1.760 ;
        RECT  1.765 0.325 2.895 0.485 ;
        RECT  2.785 0.770 2.805 1.760 ;
        RECT  2.715 0.770 2.785 1.315 ;
        RECT  2.645 0.665 2.715 1.315 ;
        RECT  2.455 0.665 2.645 0.930 ;
        RECT  2.460 2.280 2.620 2.545 ;
        RECT  2.445 1.585 2.605 2.100 ;
        RECT  1.260 2.385 2.460 2.545 ;
        RECT  2.380 1.585 2.445 1.745 ;
        RECT  2.220 1.150 2.380 1.745 ;
        RECT  1.600 2.045 2.265 2.205 ;
        RECT  2.205 1.150 2.220 1.310 ;
        RECT  2.045 0.665 2.205 1.310 ;
        RECT  1.945 0.665 2.045 0.825 ;
        RECT  1.765 1.600 2.040 1.760 ;
        RECT  1.605 0.325 1.765 1.760 ;
        RECT  1.440 1.940 1.600 2.205 ;
        RECT  1.355 1.940 1.440 2.100 ;
        RECT  1.195 0.615 1.355 2.100 ;
        RECT  1.100 2.280 1.260 2.545 ;
        RECT  0.985 2.280 1.100 2.440 ;
        RECT  0.825 0.865 0.985 2.440 ;
        RECT  0.335 0.865 0.825 1.025 ;
        RECT  0.335 2.280 0.825 2.440 ;
        RECT  0.175 0.425 0.335 1.025 ;
        RECT  0.175 2.170 0.335 2.440 ;
    END
END ADDFXLMTH

MACRO ADDHX1MTH
    CLASS CORE ;
    FOREIGN ADDHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 0.655 2.375 1.170 ;
        RECT  2.145 0.655 2.325 2.150 ;
        RECT  2.115 0.655 2.145 0.815 ;
        END
        AntennaDiffArea 0.258 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 0.765 5.230 2.005 ;
        RECT  4.945 0.765 5.020 1.025 ;
        RECT  4.945 1.745 5.020 2.005 ;
        END
        AntennaDiffArea 0.333 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.925 1.335 4.085 1.595 ;
        RECT  3.595 1.435 3.925 1.595 ;
        RECT  3.435 1.435 3.595 1.700 ;
        RECT  2.775 1.540 3.435 1.700 ;
        RECT  2.665 1.110 2.775 1.700 ;
        RECT  2.560 1.110 2.665 2.550 ;
        RECT  2.505 1.540 2.560 2.550 ;
        RECT  1.945 2.390 2.505 2.550 ;
        END
        AntennaGateArea 0.2015 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.880 3.255 1.360 ;
        END
        AntennaGateArea 0.2184 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.065 -0.130 5.330 0.130 ;
        RECT  4.125 -0.130 5.065 0.300 ;
        RECT  3.845 -0.130 4.125 0.130 ;
        RECT  3.245 -0.130 3.845 0.300 ;
        RECT  1.085 -0.130 3.245 0.130 ;
        RECT  0.145 -0.130 1.085 0.250 ;
        RECT  0.000 -0.130 0.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.645 2.740 5.330 3.000 ;
        RECT  4.385 2.570 4.645 3.000 ;
        RECT  3.595 2.740 4.385 3.000 ;
        RECT  3.335 2.570 3.595 3.000 ;
        RECT  1.280 2.740 3.335 3.000 ;
        RECT  0.340 2.620 1.280 3.000 ;
        RECT  0.000 2.740 0.340 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.765 1.220 4.790 1.480 ;
        RECT  4.605 0.655 4.765 2.380 ;
        RECT  4.015 0.655 4.605 0.815 ;
        RECT  4.105 2.220 4.605 2.380 ;
        RECT  4.265 0.995 4.425 1.935 ;
        RECT  3.595 0.995 4.265 1.155 ;
        RECT  3.935 1.775 4.265 1.935 ;
        RECT  3.845 2.220 4.105 2.420 ;
        RECT  3.775 1.775 3.935 2.040 ;
        RECT  3.005 1.880 3.775 2.040 ;
        RECT  3.435 0.480 3.595 1.155 ;
        RECT  2.785 0.480 3.435 0.640 ;
        RECT  2.845 1.880 3.005 2.360 ;
        RECT  2.625 0.310 2.785 0.640 ;
        RECT  1.425 0.310 2.625 0.470 ;
        RECT  1.765 0.655 1.905 2.120 ;
        RECT  1.745 0.655 1.765 2.410 ;
        RECT  1.605 0.655 1.745 0.815 ;
        RECT  1.605 1.960 1.745 2.410 ;
        RECT  0.385 2.250 1.605 2.410 ;
        RECT  1.355 1.180 1.565 1.440 ;
        RECT  1.265 0.310 1.425 0.635 ;
        RECT  1.195 0.815 1.355 2.070 ;
        RECT  0.755 0.475 1.265 0.635 ;
        RECT  1.095 0.815 1.195 0.975 ;
        RECT  1.095 1.910 1.195 2.070 ;
        RECT  0.595 0.475 0.755 1.540 ;
        RECT  0.465 1.280 0.595 1.540 ;
        RECT  0.285 0.735 0.385 0.995 ;
        RECT  0.285 1.995 0.385 2.410 ;
        RECT  0.125 0.735 0.285 2.410 ;
    END
END ADDHX1MTH

MACRO ADDHX2MTH
    CLASS CORE ;
    FOREIGN ADDHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.905 1.700 3.180 2.055 ;
        RECT  2.745 1.365 2.905 2.055 ;
        RECT  2.475 1.365 2.745 1.525 ;
        RECT  2.495 1.895 2.745 2.055 ;
        RECT  2.335 1.895 2.495 2.155 ;
        RECT  2.315 0.695 2.475 1.525 ;
        RECT  2.215 0.695 2.315 0.855 ;
        END
        AntennaDiffArea 0.692 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.795 1.290 6.870 1.580 ;
        RECT  6.635 0.385 6.795 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.325 1.220 3.640 1.480 ;
        RECT  3.165 0.855 3.325 1.480 ;
        RECT  2.815 0.855 3.165 1.115 ;
        RECT  2.655 0.355 2.815 1.115 ;
        RECT  1.325 0.355 2.655 0.515 ;
        RECT  1.325 1.175 1.455 1.435 ;
        RECT  1.165 0.355 1.325 1.435 ;
        RECT  0.720 1.275 1.165 1.435 ;
        RECT  0.465 1.275 0.720 1.580 ;
        END
        AntennaGateArea 0.3471 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.140 5.155 1.300 ;
        RECT  4.610 0.880 4.820 1.300 ;
        RECT  4.555 1.140 4.610 1.300 ;
        END
        AntennaGateArea 0.6006 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.305 -0.130 6.970 0.130 ;
        RECT  6.045 -0.130 6.305 0.300 ;
        RECT  4.375 -0.130 6.045 0.130 ;
        RECT  4.215 -0.130 4.375 0.300 ;
        RECT  0.825 -0.130 4.215 0.130 ;
        RECT  0.225 -0.130 0.825 0.300 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 2.740 6.970 3.000 ;
        RECT  6.075 2.205 6.335 3.000 ;
        RECT  4.425 2.740 6.075 3.000 ;
        RECT  3.485 2.620 4.425 3.000 ;
        RECT  0.820 2.740 3.485 3.000 ;
        RECT  0.220 2.465 0.820 3.000 ;
        RECT  0.000 2.740 0.220 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.225 0.820 6.385 1.855 ;
        RECT  5.905 0.820 6.225 0.980 ;
        RECT  5.935 1.695 6.225 1.855 ;
        RECT  5.495 1.225 6.045 1.485 ;
        RECT  5.675 1.695 5.935 1.980 ;
        RECT  5.645 0.720 5.905 0.980 ;
        RECT  4.975 1.820 5.675 1.980 ;
        RECT  5.320 0.720 5.645 0.880 ;
        RECT  5.335 1.225 5.495 1.640 ;
        RECT  4.015 1.480 5.335 1.640 ;
        RECT  5.160 0.540 5.320 0.880 ;
        RECT  4.035 0.540 5.160 0.700 ;
        RECT  4.875 1.820 4.975 2.200 ;
        RECT  4.715 1.820 4.875 2.440 ;
        RECT  3.055 2.280 4.715 2.440 ;
        RECT  3.875 0.310 4.035 0.700 ;
        RECT  3.855 0.880 4.015 2.005 ;
        RECT  3.155 0.310 3.875 0.470 ;
        RECT  3.665 0.880 3.855 1.040 ;
        RECT  3.815 1.745 3.855 2.005 ;
        RECT  3.505 0.650 3.665 1.040 ;
        RECT  2.995 0.310 3.155 0.615 ;
        RECT  2.795 2.280 3.055 2.560 ;
        RECT  1.365 2.400 2.795 2.560 ;
        RECT  1.975 1.125 2.135 2.220 ;
        RECT  1.065 2.060 1.975 2.220 ;
        RECT  1.635 0.695 1.795 1.875 ;
        RECT  1.505 0.695 1.635 0.855 ;
        RECT  1.245 1.715 1.635 1.875 ;
        RECT  0.905 1.805 1.065 2.220 ;
        RECT  0.385 1.805 0.905 1.965 ;
        RECT  0.285 0.745 0.385 1.005 ;
        RECT  0.285 1.755 0.385 1.965 ;
        RECT  0.125 0.745 0.285 1.965 ;
    END
END ADDHX2MTH

MACRO ADDHX4MTH
    CLASS CORE ;
    FOREIGN ADDHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.535 0.695 4.645 0.855 ;
        RECT  3.590 1.760 4.505 1.920 ;
        RECT  3.380 1.675 3.590 1.990 ;
        RECT  3.275 0.595 3.535 0.855 ;
        RECT  3.195 1.720 3.380 1.905 ;
        RECT  2.635 0.695 3.275 0.855 ;
        RECT  2.635 1.720 3.195 1.880 ;
        RECT  2.475 0.695 2.635 1.880 ;
        RECT  2.195 0.695 2.475 0.855 ;
        RECT  2.145 1.690 2.475 1.880 ;
        END
        AntennaDiffArea 1.475 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.615 1.290 9.740 1.580 ;
        RECT  9.355 0.425 9.615 2.405 ;
        END
        AntennaDiffArea 0.6 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.520 1.035 4.560 1.295 ;
        RECT  4.200 1.035 4.520 1.580 ;
        RECT  3.240 1.255 4.200 1.415 ;
        RECT  3.080 1.255 3.240 1.535 ;
        RECT  2.855 1.375 3.080 1.535 ;
        END
        AntennaGateArea 0.689 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.050 1.185 7.845 1.345 ;
        RECT  5.840 0.880 6.050 1.345 ;
        RECT  5.545 1.185 5.840 1.345 ;
        END
        AntennaGateArea 1.1973 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.125 -0.130 10.250 0.130 ;
        RECT  9.865 -0.130 10.125 0.985 ;
        RECT  9.075 -0.130 9.865 0.130 ;
        RECT  8.815 -0.130 9.075 0.590 ;
        RECT  8.025 -0.130 8.815 0.130 ;
        RECT  7.765 -0.130 8.025 0.600 ;
        RECT  6.005 -0.130 7.765 0.130 ;
        RECT  5.745 -0.130 6.005 0.300 ;
        RECT  0.385 -0.130 5.745 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.125 2.740 10.250 3.000 ;
        RECT  9.865 1.805 10.125 3.000 ;
        RECT  9.075 2.740 9.865 3.000 ;
        RECT  8.815 2.315 9.075 3.000 ;
        RECT  8.075 2.740 8.815 3.000 ;
        RECT  7.815 2.220 8.075 3.000 ;
        RECT  6.065 2.740 7.815 3.000 ;
        RECT  5.805 2.570 6.065 3.000 ;
        RECT  4.985 2.740 5.805 3.000 ;
        RECT  4.725 2.570 4.985 3.000 ;
        RECT  0.335 2.740 4.725 3.000 ;
        RECT  0.175 2.570 0.335 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.015 0.815 9.175 2.025 ;
        RECT  8.565 0.815 9.015 0.975 ;
        RECT  7.535 1.865 9.015 2.025 ;
        RECT  8.575 1.225 8.835 1.485 ;
        RECT  8.405 1.325 8.575 1.485 ;
        RECT  8.305 0.545 8.565 0.975 ;
        RECT  8.245 1.325 8.405 1.685 ;
        RECT  7.485 0.815 8.305 0.975 ;
        RECT  5.475 1.525 8.245 1.685 ;
        RECT  7.275 1.865 7.535 2.465 ;
        RECT  7.225 0.375 7.485 0.975 ;
        RECT  6.605 1.865 7.275 2.025 ;
        RECT  6.545 0.815 7.225 0.975 ;
        RECT  6.345 1.865 6.605 2.465 ;
        RECT  6.285 0.375 6.545 0.975 ;
        RECT  3.945 2.130 6.345 2.290 ;
        RECT  5.550 0.540 6.285 0.700 ;
        RECT  5.390 0.355 5.550 0.700 ;
        RECT  5.315 1.525 5.475 1.950 ;
        RECT  3.845 0.355 5.390 0.515 ;
        RECT  5.155 1.525 5.315 1.685 ;
        RECT  4.995 0.765 5.155 1.685 ;
        RECT  4.895 0.765 4.995 1.025 ;
        RECT  3.785 2.130 3.945 2.560 ;
        RECT  0.675 2.400 3.785 2.560 ;
        RECT  1.015 0.355 2.995 0.515 ;
        RECT  1.015 2.060 2.945 2.220 ;
        RECT  1.895 1.065 2.295 1.290 ;
        RECT  1.735 0.695 1.895 1.865 ;
        RECT  1.605 0.695 1.735 0.855 ;
        RECT  1.635 1.705 1.735 1.865 ;
        RECT  0.855 0.355 1.015 2.220 ;
        RECT  0.635 0.355 0.855 0.955 ;
        RECT  0.715 1.785 0.855 2.045 ;
        RECT  0.535 2.230 0.675 2.560 ;
        RECT  0.535 1.225 0.640 1.485 ;
        RECT  0.515 1.225 0.535 2.560 ;
        RECT  0.375 1.225 0.515 2.390 ;
    END
END ADDHX4MTH

MACRO ADDHX8MTH
    CLASS CORE ;
    FOREIGN ADDHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.040 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.750 0.315 8.100 1.990 ;
        RECT  7.010 0.315 7.750 0.575 ;
        RECT  6.750 0.315 7.010 2.170 ;
        RECT  5.990 0.315 6.750 0.575 ;
        RECT  5.730 0.315 5.990 2.220 ;
        RECT  4.940 2.030 5.730 2.220 ;
        RECT  4.680 0.755 4.940 2.220 ;
        RECT  3.945 2.030 4.680 2.220 ;
        RECT  3.705 0.705 3.945 2.220 ;
        END
        AntennaDiffArea 2.342 ;
    END S
    PIN CO
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.145 0.425 17.405 2.300 ;
        RECT  16.790 0.765 17.145 1.965 ;
        RECT  16.380 0.765 16.790 1.025 ;
        RECT  16.380 1.705 16.790 1.965 ;
        RECT  16.120 0.425 16.380 1.025 ;
        RECT  16.120 1.705 16.380 2.305 ;
        END
        AntennaDiffArea 1.2 ;
    END CO
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.295 1.290 3.135 1.580 ;
        END
        AntennaGateArea 1.3065 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.350 1.205 10.660 1.580 ;
        RECT  9.820 1.205 10.350 1.465 ;
        END
        AntennaGateArea 2.3881 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.915 -0.130 18.040 0.130 ;
        RECT  17.655 -0.130 17.915 1.025 ;
        RECT  16.895 -0.130 17.655 0.130 ;
        RECT  16.635 -0.130 16.895 0.565 ;
        RECT  14.910 -0.130 16.635 0.130 ;
        RECT  14.650 -0.130 14.910 0.250 ;
        RECT  11.960 -0.130 14.650 0.130 ;
        RECT  11.700 -0.130 11.960 0.250 ;
        RECT  9.930 -0.130 11.700 0.130 ;
        RECT  9.670 -0.130 9.930 0.250 ;
        RECT  3.175 -0.130 9.670 0.130 ;
        RECT  2.915 -0.130 3.175 0.250 ;
        RECT  0.385 -0.130 2.915 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.915 2.740 18.040 3.000 ;
        RECT  17.655 1.785 17.915 3.000 ;
        RECT  16.895 2.740 17.655 3.000 ;
        RECT  16.635 2.155 16.895 3.000 ;
        RECT  15.870 2.740 16.635 3.000 ;
        RECT  15.610 1.895 15.870 3.000 ;
        RECT  14.850 2.740 15.610 3.000 ;
        RECT  14.590 1.895 14.850 3.000 ;
        RECT  13.830 2.740 14.590 3.000 ;
        RECT  13.570 1.895 13.830 3.000 ;
        RECT  12.810 2.740 13.570 3.000 ;
        RECT  12.550 1.895 12.810 3.000 ;
        RECT  11.790 2.740 12.550 3.000 ;
        RECT  11.530 1.895 11.790 3.000 ;
        RECT  10.740 2.740 11.530 3.000 ;
        RECT  10.480 2.570 10.740 3.000 ;
        RECT  9.660 2.740 10.480 3.000 ;
        RECT  9.400 2.570 9.660 3.000 ;
        RECT  8.560 2.740 9.400 3.000 ;
        RECT  8.300 2.570 8.560 3.000 ;
        RECT  3.155 2.740 8.300 3.000 ;
        RECT  2.215 2.620 3.155 3.000 ;
        RECT  0.385 2.740 2.215 3.000 ;
        RECT  0.125 2.465 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.885 1.265 16.565 1.525 ;
        RECT  15.725 0.445 15.885 1.525 ;
        RECT  10.850 0.445 15.725 0.605 ;
        RECT  15.360 0.785 15.450 1.385 ;
        RECT  15.190 0.785 15.360 2.285 ;
        RECT  15.100 1.185 15.190 2.285 ;
        RECT  14.370 1.185 15.100 1.385 ;
        RECT  14.340 0.785 14.370 1.385 ;
        RECT  14.110 0.785 14.340 2.285 ;
        RECT  14.080 1.185 14.110 2.285 ;
        RECT  13.430 1.185 14.080 1.385 ;
        RECT  13.320 0.785 13.430 1.385 ;
        RECT  13.170 0.785 13.320 2.285 ;
        RECT  13.060 1.185 13.170 2.285 ;
        RECT  12.500 1.185 13.060 1.385 ;
        RECT  12.300 0.785 12.500 1.385 ;
        RECT  12.240 0.785 12.300 2.285 ;
        RECT  12.040 1.185 12.240 2.285 ;
        RECT  11.410 1.185 12.040 1.385 ;
        RECT  11.280 0.785 11.410 1.385 ;
        RECT  11.150 0.785 11.280 2.380 ;
        RECT  11.020 1.185 11.150 2.380 ;
        RECT  7.490 2.220 11.020 2.380 ;
        RECT  10.690 0.445 10.850 0.975 ;
        RECT  8.920 0.815 10.690 0.975 ;
        RECT  10.210 0.355 10.470 0.635 ;
        RECT  9.020 0.475 10.210 0.635 ;
        RECT  9.940 1.770 10.200 2.030 ;
        RECT  9.120 1.870 9.940 2.030 ;
        RECT  8.920 1.770 9.120 2.030 ;
        RECT  8.760 0.355 9.020 0.635 ;
        RECT  8.760 0.815 8.920 2.030 ;
        RECT  8.510 0.815 8.760 0.975 ;
        RECT  8.280 0.375 8.510 0.975 ;
        RECT  7.230 0.755 7.490 2.560 ;
        RECT  6.470 2.400 7.230 2.560 ;
        RECT  6.210 0.755 6.470 2.560 ;
        RECT  3.495 2.400 6.210 2.560 ;
        RECT  5.220 0.365 5.480 1.850 ;
        RECT  4.455 0.365 5.220 0.525 ;
        RECT  4.195 0.365 4.455 1.850 ;
        RECT  3.515 0.365 4.195 0.525 ;
        RECT  3.365 0.835 3.525 2.100 ;
        RECT  3.355 0.365 3.515 0.635 ;
        RECT  3.335 2.280 3.495 2.560 ;
        RECT  3.335 0.835 3.365 1.095 ;
        RECT  2.545 1.785 3.365 1.945 ;
        RECT  1.855 0.475 3.355 0.635 ;
        RECT  2.775 0.890 3.335 1.050 ;
        RECT  3.095 2.280 3.335 2.440 ;
        RECT  2.935 2.125 3.095 2.440 ;
        RECT  0.485 2.125 2.935 2.285 ;
        RECT  2.515 0.815 2.775 1.050 ;
        RECT  1.825 0.330 1.855 0.635 ;
        RECT  1.825 0.830 1.855 1.895 ;
        RECT  1.595 0.330 1.825 1.895 ;
        RECT  1.565 0.330 1.595 1.025 ;
        RECT  0.665 1.735 1.595 1.895 ;
        RECT  0.895 0.330 1.565 0.490 ;
        RECT  0.485 1.225 1.315 1.485 ;
        RECT  0.635 0.330 0.895 1.025 ;
        RECT  0.325 1.225 0.485 2.285 ;
    END
END ADDHX8MTH

MACRO AND2X12MTH
    CLASS CORE ;
    FOREIGN AND2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.705 1.725 2.965 2.410 ;
        RECT  2.645 0.385 2.905 1.105 ;
        RECT  1.945 1.725 2.705 2.095 ;
        RECT  1.945 0.745 2.645 1.105 ;
        RECT  1.685 0.385 1.945 2.410 ;
        RECT  1.620 0.385 1.685 1.785 ;
        RECT  0.925 1.085 1.620 1.785 ;
        RECT  0.665 0.385 0.925 2.410 ;
        END
        AntennaDiffArea 1.806 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.560 1.250 4.500 1.580 ;
        END
        AntennaGateArea 0.4641 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.965 1.230 5.585 1.580 ;
        END
        AntennaGateArea 0.4641 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 -0.130 6.560 0.130 ;
        RECT  4.120 -0.130 4.380 0.685 ;
        RECT  2.390 -0.130 4.120 0.130 ;
        RECT  2.130 -0.130 2.390 0.565 ;
        RECT  0.385 -0.130 2.130 0.130 ;
        RECT  0.125 -0.130 0.385 0.995 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.885 6.435 3.000 ;
        RECT  4.435 2.740 6.175 3.000 ;
        RECT  4.175 2.140 4.435 3.000 ;
        RECT  2.455 2.740 4.175 3.000 ;
        RECT  2.195 2.275 2.455 3.000 ;
        RECT  1.435 2.740 2.195 3.000 ;
        RECT  1.175 2.180 1.435 3.000 ;
        RECT  0.385 2.740 1.175 3.000 ;
        RECT  0.125 2.025 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.175 0.765 6.435 1.040 ;
        RECT  5.925 0.880 6.175 1.040 ;
        RECT  5.665 0.455 5.925 0.685 ;
        RECT  5.890 0.880 5.925 1.960 ;
        RECT  5.765 0.880 5.890 2.160 ;
        RECT  5.415 0.880 5.765 1.040 ;
        RECT  5.630 1.800 5.765 2.160 ;
        RECT  4.900 0.455 5.665 0.615 ;
        RECT  4.955 1.800 5.630 1.960 ;
        RECT  5.155 0.815 5.415 1.040 ;
        RECT  4.695 1.800 4.955 2.275 ;
        RECT  4.740 0.455 4.900 1.025 ;
        RECT  4.640 0.750 4.740 1.025 ;
        RECT  3.915 1.800 4.695 1.960 ;
        RECT  3.860 0.865 4.640 1.025 ;
        RECT  3.655 1.800 3.915 2.275 ;
        RECT  3.600 0.765 3.860 1.025 ;
        RECT  3.305 1.800 3.655 1.960 ;
        RECT  3.145 1.285 3.305 1.960 ;
        RECT  2.195 1.285 3.145 1.545 ;
    END
END AND2X12MTH

MACRO AND2X1MTH
    CLASS CORE ;
    FOREIGN AND2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.880 0.715 1.950 1.235 ;
        RECT  1.690 0.715 1.880 2.280 ;
        END
        AntennaDiffArea 0.329 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.290 1.170 1.780 ;
        END
        AntennaGateArea 0.0598 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.285 0.580 1.635 ;
        END
        AntennaGateArea 0.0598 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 -0.130 2.050 0.130 ;
        RECT  1.665 -0.130 1.925 0.300 ;
        RECT  1.385 -0.130 1.665 0.130 ;
        RECT  0.445 -0.130 1.385 0.300 ;
        RECT  0.000 -0.130 0.445 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.385 2.740 2.050 3.000 ;
        RECT  1.125 2.570 1.385 3.000 ;
        RECT  0.725 2.740 1.125 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.350 0.885 1.510 2.150 ;
        RECT  0.385 0.885 1.350 1.045 ;
        RECT  0.635 1.990 1.350 2.150 ;
        RECT  0.125 0.765 0.385 1.045 ;
    END
END AND2X1MTH

MACRO AND2X2MTH
    CLASS CORE ;
    FOREIGN AND2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 0.470 1.950 0.760 ;
        RECT  1.695 0.470 1.875 2.405 ;
        RECT  1.665 0.470 1.695 0.760 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.755 1.290 1.165 1.760 ;
        END
        AntennaGateArea 0.0962 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.285 0.470 1.735 ;
        END
        AntennaGateArea 0.0962 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.130 2.050 0.130 ;
        RECT  1.050 -0.130 1.310 0.640 ;
        RECT  0.750 -0.130 1.050 0.130 ;
        RECT  0.150 -0.130 0.750 0.300 ;
        RECT  0.000 -0.130 0.150 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.385 2.740 2.050 3.000 ;
        RECT  1.125 2.280 1.385 3.000 ;
        RECT  0.785 2.570 1.125 3.000 ;
        RECT  0.385 2.740 0.785 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.350 0.885 1.510 2.100 ;
        RECT  0.385 0.885 1.350 1.045 ;
        RECT  0.835 1.940 1.350 2.100 ;
        RECT  0.575 1.940 0.835 2.270 ;
        RECT  0.125 0.745 0.385 1.045 ;
    END
END AND2X2MTH

MACRO AND2X4MTH
    CLASS CORE ;
    FOREIGN AND2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.715 1.270 2.770 1.605 ;
        RECT  2.535 0.390 2.715 2.420 ;
        RECT  2.405 0.390 2.535 0.990 ;
        RECT  2.425 1.820 2.535 2.420 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 0.950 1.815 1.840 ;
        RECT  0.485 0.950 1.655 1.110 ;
        RECT  0.325 0.870 0.485 1.750 ;
        RECT  0.100 0.870 0.325 1.170 ;
        END
        AntennaGateArea 0.1924 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.780 1.290 1.190 1.745 ;
        END
        AntennaGateArea 0.1924 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 -0.130 3.280 0.130 ;
        RECT  2.895 -0.130 3.155 0.980 ;
        RECT  2.075 -0.130 2.895 0.130 ;
        RECT  1.815 -0.130 2.075 0.300 ;
        RECT  0.725 -0.130 1.815 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 2.740 3.280 3.000 ;
        RECT  1.870 2.570 2.130 3.000 ;
        RECT  1.580 2.740 1.870 3.000 ;
        RECT  0.980 2.570 1.580 3.000 ;
        RECT  0.725 2.740 0.980 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.225 1.145 2.290 1.405 ;
        RECT  2.065 0.610 2.225 2.215 ;
        RECT  0.955 0.610 2.065 0.770 ;
        RECT  0.510 2.055 2.065 2.215 ;
    END
END AND2X4MTH

MACRO AND2X6MTH
    CLASS CORE ;
    FOREIGN AND2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.705 0.390 3.975 2.420 ;
        RECT  2.955 1.280 3.705 1.580 ;
        RECT  2.685 0.385 2.955 2.420 ;
        END
        AntennaDiffArea 1.169 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.285 1.985 1.545 ;
        RECT  1.725 0.955 1.885 1.545 ;
        RECT  0.720 0.955 1.725 1.115 ;
        RECT  0.595 0.880 0.720 1.170 ;
        RECT  0.335 0.880 0.595 1.565 ;
        END
        AntennaGateArea 0.234 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.330 1.480 1.655 ;
        END
        AntennaGateArea 0.234 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 -0.130 4.100 0.130 ;
        RECT  3.175 -0.130 3.435 1.005 ;
        RECT  2.250 -0.130 3.175 0.130 ;
        RECT  1.990 -0.130 2.250 0.300 ;
        RECT  1.450 -0.130 1.990 0.130 ;
        RECT  0.850 -0.130 1.450 0.300 ;
        RECT  0.385 -0.130 0.850 0.130 ;
        RECT  0.125 -0.130 0.385 0.670 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  3.175 1.820 3.435 3.000 ;
        RECT  2.355 2.740 3.175 3.000 ;
        RECT  2.095 2.230 2.355 3.000 ;
        RECT  1.685 2.740 2.095 3.000 ;
        RECT  1.085 2.570 1.685 3.000 ;
        RECT  0.725 2.740 1.085 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.345 1.220 2.505 1.480 ;
        RECT  2.185 0.615 2.345 1.995 ;
        RECT  1.015 0.615 2.185 0.775 ;
        RECT  1.800 1.835 2.185 1.995 ;
        RECT  1.540 1.835 1.800 2.095 ;
        RECT  0.805 1.835 1.540 1.995 ;
        RECT  0.545 1.835 0.805 2.095 ;
    END
END AND2X6MTH

MACRO AND2X8MTH
    CLASS CORE ;
    FOREIGN AND2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.580 0.390 3.840 2.440 ;
        RECT  3.375 0.640 3.580 1.970 ;
        RECT  2.760 0.640 3.375 0.990 ;
        RECT  2.760 1.620 3.375 1.970 ;
        RECT  2.500 0.390 2.760 0.990 ;
        RECT  2.500 1.620 2.760 2.440 ;
        END
        AntennaDiffArea 1.208 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.805 1.240 1.965 1.795 ;
        RECT  0.720 1.635 1.805 1.795 ;
        RECT  0.405 1.245 0.720 1.795 ;
        END
        AntennaGateArea 0.3094 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 0.880 1.550 1.455 ;
        END
        AntennaGateArea 0.3094 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  4.125 -0.130 4.385 0.980 ;
        RECT  3.300 -0.130 4.125 0.130 ;
        RECT  3.040 -0.130 3.300 0.455 ;
        RECT  2.220 -0.130 3.040 0.130 ;
        RECT  1.960 -0.130 2.220 0.300 ;
        RECT  0.405 -0.130 1.960 0.130 ;
        RECT  0.145 -0.130 0.405 0.980 ;
        RECT  0.000 -0.130 0.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.755 4.385 3.000 ;
        RECT  3.300 2.740 4.125 3.000 ;
        RECT  3.040 2.155 3.300 3.000 ;
        RECT  2.220 2.740 3.040 3.000 ;
        RECT  1.620 2.570 2.220 3.000 ;
        RECT  1.310 2.740 1.620 3.000 ;
        RECT  1.050 2.570 1.310 3.000 ;
        RECT  0.725 2.740 1.050 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.305 1.175 2.930 1.435 ;
        RECT  2.145 0.525 2.305 2.140 ;
        RECT  1.075 0.525 2.145 0.685 ;
        RECT  1.725 1.980 2.145 2.140 ;
        RECT  1.465 1.980 1.725 2.240 ;
        RECT  0.795 1.980 1.465 2.140 ;
        RECT  0.535 1.980 0.795 2.240 ;
    END
END AND2X8MTH

MACRO AND3X12MTH
    CLASS CORE ;
    FOREIGN AND3X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.635 0.385 2.855 0.985 ;
        RECT  2.635 1.810 2.785 2.410 ;
        RECT  2.335 0.385 2.635 2.410 ;
        RECT  1.935 1.085 2.335 1.785 ;
        RECT  1.855 0.385 1.935 1.785 ;
        RECT  1.675 0.385 1.855 2.410 ;
        RECT  1.595 1.085 1.675 2.410 ;
        RECT  0.925 1.085 1.595 1.785 ;
        RECT  0.665 0.385 0.925 2.410 ;
        END
        AntennaDiffArea 1.8 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 1.125 6.345 1.345 ;
        RECT  5.675 0.770 5.835 1.345 ;
        RECT  3.715 0.770 5.675 0.930 ;
        RECT  3.555 0.770 3.715 1.580 ;
        RECT  3.375 1.230 3.555 1.580 ;
        END
        AntennaGateArea 0.507 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.585 2.240 6.845 2.555 ;
        RECT  5.545 2.240 6.585 2.400 ;
        RECT  5.285 2.240 5.545 2.555 ;
        RECT  4.040 2.240 5.285 2.400 ;
        RECT  3.905 2.140 4.040 2.400 ;
        RECT  3.645 2.140 3.905 2.560 ;
        END
        AntennaGateArea 0.507 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.030 1.230 7.385 1.685 ;
        RECT  5.095 1.525 7.030 1.685 ;
        RECT  4.935 1.230 5.095 1.685 ;
        RECT  4.325 1.230 4.935 1.490 ;
        END
        AntennaGateArea 0.507 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.170 -0.130 7.790 0.130 ;
        RECT  5.910 -0.130 6.170 0.250 ;
        RECT  3.495 -0.130 5.910 0.130 ;
        RECT  3.235 -0.130 3.495 0.250 ;
        RECT  0.385 -0.130 3.235 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.625 2.740 7.790 3.000 ;
        RECT  7.025 2.570 7.625 3.000 ;
        RECT  6.405 2.740 7.025 3.000 ;
        RECT  5.805 2.620 6.405 3.000 ;
        RECT  5.115 2.740 5.805 3.000 ;
        RECT  4.855 2.620 5.115 3.000 ;
        RECT  4.675 2.740 4.855 3.000 ;
        RECT  4.075 2.620 4.675 3.000 ;
        RECT  3.325 2.740 4.075 3.000 ;
        RECT  3.065 2.570 3.325 3.000 ;
        RECT  0.385 2.740 3.065 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.405 1.880 7.665 2.140 ;
        RECT  7.235 0.390 7.495 0.990 ;
        RECT  4.735 1.880 7.405 2.040 ;
        RECT  3.195 0.430 7.235 0.590 ;
        RECT  4.475 1.780 4.735 2.040 ;
        RECT  3.195 1.780 4.475 1.940 ;
        RECT  3.035 0.430 3.195 1.940 ;
        RECT  2.815 1.235 3.035 1.495 ;
    END
END AND3X12MTH

MACRO AND3X1MTH
    CLASS CORE ;
    FOREIGN AND3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 0.760 2.360 1.170 ;
        RECT  2.175 0.760 2.335 2.010 ;
        RECT  2.150 0.760 2.175 1.170 ;
        RECT  2.125 1.750 2.175 2.010 ;
        RECT  2.075 0.760 2.150 1.020 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 0.880 1.540 1.515 ;
        END
        AntennaGateArea 0.0663 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.460 1.130 1.235 ;
        RECT  0.825 0.460 0.900 0.620 ;
        END
        AntennaGateArea 0.0663 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.220 0.720 1.795 ;
        END
        AntennaGateArea 0.0663 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 -0.130 2.460 0.130 ;
        RECT  1.790 -0.130 2.130 0.300 ;
        RECT  1.530 -0.130 1.790 0.645 ;
        RECT  1.110 -0.130 1.530 0.130 ;
        RECT  0.170 -0.130 1.110 0.250 ;
        RECT  0.000 -0.130 0.170 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.275 2.740 2.460 3.000 ;
        RECT  1.675 2.555 2.275 3.000 ;
        RECT  0.895 2.740 1.675 3.000 ;
        RECT  0.635 2.445 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.935 1.295 1.995 1.555 ;
        RECT  1.775 1.295 1.935 2.235 ;
        RECT  1.405 2.075 1.775 2.235 ;
        RECT  1.145 2.075 1.405 2.445 ;
        RECT  0.385 2.075 1.145 2.235 ;
        RECT  0.285 0.760 0.385 1.020 ;
        RECT  0.285 2.075 0.385 2.430 ;
        RECT  0.125 0.760 0.285 2.430 ;
    END
END AND3X1MTH

MACRO AND3X2MTH
    CLASS CORE ;
    FOREIGN AND3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 0.385 2.365 2.355 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 1.055 1.540 1.580 ;
        END
        AntennaGateArea 0.1066 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.035 1.700 1.130 1.990 ;
        RECT  0.775 1.255 1.035 1.990 ;
        END
        AntennaGateArea 0.1066 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.260 0.555 1.600 ;
        END
        AntennaGateArea 0.1066 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.795 -0.130 2.460 0.130 ;
        RECT  1.195 -0.130 1.795 0.300 ;
        RECT  0.785 -0.130 1.195 0.130 ;
        RECT  0.185 -0.130 0.785 0.300 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.795 2.740 2.460 3.000 ;
        RECT  1.535 2.620 1.795 3.000 ;
        RECT  0.775 2.740 1.535 3.000 ;
        RECT  0.175 2.620 0.775 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.785 0.665 1.945 2.440 ;
        RECT  0.385 0.665 1.785 0.825 ;
        RECT  1.285 2.280 1.785 2.440 ;
        RECT  1.025 2.280 1.285 2.515 ;
        RECT  0.385 2.280 1.025 2.440 ;
        RECT  0.125 0.665 0.385 0.925 ;
        RECT  0.125 1.780 0.385 2.440 ;
    END
END AND3X2MTH

MACRO AND3X4MTH
    CLASS CORE ;
    FOREIGN AND3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.235 2.770 1.595 ;
        RECT  2.295 1.235 2.335 2.310 ;
        RECT  2.135 0.445 2.295 2.310 ;
        RECT  1.945 0.445 2.135 0.605 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.135 1.570 1.605 ;
        END
        AntennaGateArea 0.1885 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.790 1.135 1.130 1.605 ;
        END
        AntennaGateArea 0.1885 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.165 0.510 1.605 ;
        END
        AntennaGateArea 0.1885 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 2.870 0.130 ;
        RECT  2.485 -0.130 2.745 1.000 ;
        RECT  1.695 -0.130 2.485 0.130 ;
        RECT  1.435 -0.130 1.695 0.615 ;
        RECT  0.000 -0.130 1.435 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.835 2.740 2.870 3.000 ;
        RECT  1.575 2.125 1.835 3.000 ;
        RECT  0.000 2.740 1.575 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.910 1.205 1.955 1.465 ;
        RECT  1.750 0.795 1.910 1.945 ;
        RECT  0.385 0.795 1.750 0.955 ;
        RECT  1.325 1.785 1.750 1.945 ;
        RECT  1.065 1.785 1.325 2.090 ;
        RECT  0.385 1.785 1.065 1.945 ;
        RECT  0.125 0.355 0.385 0.955 ;
        RECT  0.125 1.785 0.385 2.095 ;
    END
END AND3X4MTH

MACRO AND3X6MTH
    CLASS CORE ;
    FOREIGN AND3X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 0.385 5.205 2.410 ;
        RECT  4.185 1.285 4.945 1.585 ;
        RECT  3.925 0.385 4.185 2.415 ;
        RECT  3.865 0.385 3.925 0.985 ;
        END
        AntennaDiffArea 1.137 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.165 1.230 3.265 1.490 ;
        RECT  3.005 0.925 3.165 1.490 ;
        RECT  0.720 0.925 3.005 1.085 ;
        RECT  0.560 0.925 0.720 1.585 ;
        RECT  0.305 1.185 0.560 1.585 ;
        END
        AntennaGateArea 0.3224 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.275 2.675 1.585 ;
        END
        AntennaGateArea 0.3224 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.275 1.940 1.585 ;
        END
        AntennaGateArea 0.3224 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.665 -0.130 5.330 0.130 ;
        RECT  4.405 -0.130 4.665 0.990 ;
        RECT  3.475 -0.130 4.405 0.130 ;
        RECT  3.215 -0.130 3.475 0.300 ;
        RECT  0.755 -0.130 3.215 0.130 ;
        RECT  0.155 -0.130 0.755 0.640 ;
        RECT  0.000 -0.130 0.155 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.695 2.740 5.330 3.000 ;
        RECT  4.435 1.810 4.695 3.000 ;
        RECT  3.635 2.740 4.435 3.000 ;
        RECT  3.375 2.110 3.635 3.000 ;
        RECT  3.035 2.570 3.375 3.000 ;
        RECT  2.535 2.740 3.035 3.000 ;
        RECT  2.275 2.110 2.535 3.000 ;
        RECT  1.455 2.740 2.275 3.000 ;
        RECT  1.195 2.110 1.455 3.000 ;
        RECT  0.725 2.740 1.195 3.000 ;
        RECT  0.385 2.570 0.725 3.000 ;
        RECT  0.125 1.830 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.605 1.230 3.695 1.490 ;
        RECT  3.445 0.585 3.605 1.930 ;
        RECT  1.965 0.585 3.445 0.745 ;
        RECT  0.645 1.770 3.445 1.930 ;
        RECT  1.705 0.485 1.965 0.745 ;
    END
END AND3X6MTH

MACRO AND3X8MTH
    CLASS CORE ;
    FOREIGN AND3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 0.385 2.015 0.985 ;
        RECT  1.645 0.385 1.935 2.410 ;
        RECT  0.935 1.240 1.645 1.590 ;
        RECT  0.905 0.385 0.935 1.590 ;
        RECT  0.675 0.385 0.905 2.410 ;
        RECT  0.645 1.085 0.675 2.410 ;
        RECT  0.510 1.085 0.645 1.785 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.925 1.125 5.435 1.345 ;
        RECT  4.765 0.770 4.925 1.345 ;
        RECT  2.880 0.770 4.765 0.930 ;
        RECT  2.720 0.770 2.880 1.580 ;
        RECT  2.560 1.135 2.720 1.580 ;
        END
        AntennaGateArea 0.4251 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 2.245 6.020 2.455 ;
        RECT  4.710 2.245 5.760 2.405 ;
        RECT  4.450 2.245 4.710 2.455 ;
        RECT  3.220 2.245 4.450 2.405 ;
        RECT  3.165 2.140 3.220 2.405 ;
        RECT  2.900 2.140 3.165 2.455 ;
        END
        AntennaGateArea 0.4251 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.210 1.230 6.565 1.685 ;
        RECT  4.275 1.525 6.210 1.685 ;
        RECT  4.115 1.230 4.275 1.685 ;
        RECT  3.505 1.230 4.115 1.490 ;
        END
        AntennaGateArea 0.4251 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.350 -0.130 6.970 0.130 ;
        RECT  5.090 -0.130 5.350 0.250 ;
        RECT  2.595 -0.130 5.090 0.130 ;
        RECT  2.335 -0.130 2.595 0.250 ;
        RECT  1.465 -0.130 2.335 0.130 ;
        RECT  1.225 -0.130 1.465 1.000 ;
        RECT  0.395 -0.130 1.225 0.130 ;
        RECT  0.135 -0.130 0.395 0.945 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.770 2.740 6.970 3.000 ;
        RECT  6.170 2.570 6.770 3.000 ;
        RECT  5.605 2.740 6.170 3.000 ;
        RECT  5.005 2.620 5.605 3.000 ;
        RECT  4.335 2.740 5.005 3.000 ;
        RECT  4.075 2.620 4.335 3.000 ;
        RECT  3.875 2.740 4.075 3.000 ;
        RECT  3.275 2.620 3.875 3.000 ;
        RECT  2.465 2.740 3.275 3.000 ;
        RECT  2.175 2.135 2.465 3.000 ;
        RECT  1.415 2.740 2.175 3.000 ;
        RECT  1.155 1.810 1.415 3.000 ;
        RECT  0.385 2.740 1.155 3.000 ;
        RECT  0.125 1.915 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.585 1.865 6.845 2.125 ;
        RECT  6.375 0.620 6.675 0.880 ;
        RECT  3.935 1.865 6.585 2.025 ;
        RECT  6.215 0.430 6.375 0.880 ;
        RECT  2.380 0.430 6.215 0.590 ;
        RECT  3.655 1.780 3.935 2.025 ;
        RECT  2.380 1.780 3.655 1.940 ;
        RECT  2.220 0.430 2.380 1.940 ;
        RECT  2.115 1.235 2.220 1.495 ;
    END
END AND3X8MTH

MACRO AND3XLMTH
    CLASS CORE ;
    FOREIGN AND3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.760 2.360 1.945 ;
        RECT  2.150 0.760 2.200 1.170 ;
        RECT  2.125 1.685 2.200 1.945 ;
        RECT  2.075 0.760 2.150 1.020 ;
        END
        AntennaDiffArea 0.231 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 0.880 1.540 1.515 ;
        END
        AntennaGateArea 0.0533 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.500 1.130 1.235 ;
        RECT  0.825 0.500 0.900 0.760 ;
        END
        AntennaGateArea 0.0533 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.220 0.720 1.795 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 -0.130 2.460 0.130 ;
        RECT  1.530 -0.130 2.130 0.510 ;
        RECT  1.120 -0.130 1.530 0.130 ;
        RECT  0.180 -0.130 1.120 0.300 ;
        RECT  0.000 -0.130 0.180 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.275 2.740 2.460 3.000 ;
        RECT  1.675 2.460 2.275 3.000 ;
        RECT  0.895 2.740 1.675 3.000 ;
        RECT  0.635 2.560 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.935 1.295 1.995 1.555 ;
        RECT  1.775 1.295 1.935 2.235 ;
        RECT  1.405 2.075 1.775 2.235 ;
        RECT  1.145 2.075 1.405 2.425 ;
        RECT  0.385 2.075 1.145 2.235 ;
        RECT  0.285 0.760 0.385 1.020 ;
        RECT  0.285 2.075 0.385 2.430 ;
        RECT  0.125 0.760 0.285 2.430 ;
    END
END AND3XLMTH

MACRO AND4X12MTH
    CLASS CORE ;
    FOREIGN AND4X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.725 0.385 3.095 2.410 ;
        RECT  2.675 0.385 2.725 1.635 ;
        RECT  2.005 1.095 2.675 1.635 ;
        RECT  1.855 1.095 2.005 2.410 ;
        RECT  1.745 0.385 1.855 2.410 ;
        RECT  1.595 0.385 1.745 1.785 ;
        RECT  0.925 1.085 1.595 1.785 ;
        RECT  0.665 0.385 0.925 2.410 ;
        END
        AntennaDiffArea 1.8 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.010 1.280 5.290 1.560 ;
        END
        AntennaGateArea 0.6292 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.055 1.280 7.335 1.560 ;
        END
        AntennaGateArea 0.6292 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.690 1.280 9.970 1.555 ;
        END
        AntennaGateArea 0.6292 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.575 1.280 11.855 1.555 ;
        END
        AntennaGateArea 0.6292 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.300 -0.130 12.710 0.130 ;
        RECT  5.040 -0.130 5.300 0.615 ;
        RECT  2.395 -0.130 5.040 0.130 ;
        RECT  2.135 -0.130 2.395 0.640 ;
        RECT  0.385 -0.130 2.135 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.580 2.740 12.710 3.000 ;
        RECT  12.320 2.230 12.580 3.000 ;
        RECT  12.025 2.740 12.320 3.000 ;
        RECT  11.765 2.570 12.025 3.000 ;
        RECT  11.485 2.740 11.765 3.000 ;
        RECT  11.225 2.230 11.485 3.000 ;
        RECT  10.930 2.740 11.225 3.000 ;
        RECT  10.670 2.570 10.930 3.000 ;
        RECT  10.385 2.740 10.670 3.000 ;
        RECT  10.125 2.230 10.385 3.000 ;
        RECT  9.830 2.740 10.125 3.000 ;
        RECT  9.570 2.570 9.830 3.000 ;
        RECT  9.285 2.740 9.570 3.000 ;
        RECT  9.025 2.230 9.285 3.000 ;
        RECT  8.715 2.740 9.025 3.000 ;
        RECT  8.455 2.570 8.715 3.000 ;
        RECT  8.115 2.740 8.455 3.000 ;
        RECT  7.855 2.230 8.115 3.000 ;
        RECT  7.545 2.740 7.855 3.000 ;
        RECT  7.285 2.570 7.545 3.000 ;
        RECT  6.945 2.740 7.285 3.000 ;
        RECT  6.685 2.230 6.945 3.000 ;
        RECT  6.390 2.740 6.685 3.000 ;
        RECT  6.130 2.570 6.390 3.000 ;
        RECT  5.845 2.740 6.130 3.000 ;
        RECT  5.585 2.230 5.845 3.000 ;
        RECT  5.290 2.740 5.585 3.000 ;
        RECT  5.030 2.570 5.290 3.000 ;
        RECT  4.745 2.740 5.030 3.000 ;
        RECT  4.485 2.230 4.745 3.000 ;
        RECT  4.200 2.740 4.485 3.000 ;
        RECT  3.940 2.570 4.200 3.000 ;
        RECT  3.645 2.740 3.940 3.000 ;
        RECT  3.365 2.230 3.645 3.000 ;
        RECT  2.545 2.740 3.365 3.000 ;
        RECT  2.285 1.890 2.545 3.000 ;
        RECT  1.465 2.740 2.285 3.000 ;
        RECT  1.205 2.095 1.465 3.000 ;
        RECT  0.385 2.740 1.205 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.505 0.405 12.585 0.565 ;
        RECT  12.075 0.815 12.235 1.935 ;
        RECT  10.770 0.815 12.075 0.975 ;
        RECT  3.535 1.775 12.075 1.935 ;
        RECT  10.345 0.405 10.505 0.970 ;
        RECT  8.170 0.810 10.345 0.970 ;
        RECT  6.095 0.405 9.985 0.565 ;
        RECT  5.785 0.805 7.910 0.965 ;
        RECT  5.625 0.355 5.785 0.965 ;
        RECT  4.740 0.805 5.625 0.965 ;
        RECT  4.580 0.355 4.740 0.965 ;
        RECT  3.850 0.805 4.580 0.965 ;
        RECT  3.590 0.355 3.850 0.965 ;
        RECT  3.375 1.235 3.535 1.935 ;
        RECT  3.275 1.235 3.375 1.495 ;
    END
END AND4X12MTH

MACRO AND4X1MTH
    CLASS CORE ;
    FOREIGN AND4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.735 2.770 2.220 ;
        RECT  2.485 0.735 2.610 1.170 ;
        RECT  2.485 1.960 2.610 2.220 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 0.825 2.000 1.440 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 0.415 1.540 0.760 ;
        END
        AntennaGateArea 0.0728 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.805 1.300 1.150 1.990 ;
        END
        AntennaGateArea 0.0728 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.535 1.585 ;
        END
        AntennaGateArea 0.0728 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 -0.130 2.870 0.130 ;
        RECT  1.910 -0.130 2.510 0.415 ;
        RECT  0.730 -0.130 1.910 0.130 ;
        RECT  0.130 -0.130 0.730 0.300 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.190 2.740 2.870 3.000 ;
        RECT  1.590 2.620 2.190 3.000 ;
        RECT  1.320 2.740 1.590 3.000 ;
        RECT  1.060 2.620 1.320 3.000 ;
        RECT  0.000 2.740 1.060 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.180 1.380 2.400 1.780 ;
        RECT  1.760 1.620 2.180 1.780 ;
        RECT  1.520 1.620 1.760 2.400 ;
        RECT  1.500 0.940 1.520 2.400 ;
        RECT  1.360 0.940 1.500 1.780 ;
        RECT  0.810 2.240 1.500 2.400 ;
        RECT  0.385 0.940 1.360 1.100 ;
        RECT  0.550 2.240 0.810 2.500 ;
        RECT  0.125 0.765 0.385 1.100 ;
    END
END AND4X1MTH

MACRO AND4X2MTH
    CLASS CORE ;
    FOREIGN AND4X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.460 2.770 2.415 ;
        RECT  2.560 0.460 2.610 1.180 ;
        RECT  2.485 1.815 2.610 2.415 ;
        RECT  2.485 0.460 2.560 0.760 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.650 1.160 1.950 1.580 ;
        END
        AntennaGateArea 0.1183 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 2.110 1.725 2.390 ;
        END
        AntennaGateArea 0.1183 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.765 0.880 1.130 1.575 ;
        END
        AntennaGateArea 0.1183 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.340 0.965 0.395 1.225 ;
        RECT  0.100 0.965 0.340 1.590 ;
        END
        AntennaGateArea 0.1183 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.155 -0.130 2.870 0.130 ;
        RECT  1.895 -0.130 2.155 0.980 ;
        RECT  0.000 -0.130 1.895 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 2.740 2.870 3.000 ;
        RECT  1.605 2.570 2.205 3.000 ;
        RECT  1.275 2.740 1.605 3.000 ;
        RECT  1.015 2.570 1.275 3.000 ;
        RECT  0.725 2.740 1.015 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.290 1.315 2.355 1.575 ;
        RECT  2.130 1.315 2.290 1.920 ;
        RECT  1.470 1.760 2.130 1.920 ;
        RECT  1.310 0.535 1.470 1.920 ;
        RECT  0.555 0.535 1.310 0.695 ;
        RECT  0.525 1.760 1.310 1.920 ;
        RECT  0.295 0.435 0.555 0.695 ;
    END
END AND4X2MTH

MACRO AND4X4MTH
    CLASS CORE ;
    FOREIGN AND4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.665 1.245 4.860 1.580 ;
        RECT  4.485 0.395 4.665 2.415 ;
        RECT  4.455 0.395 4.485 0.995 ;
        RECT  4.455 1.815 4.485 2.415 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.340 0.770 3.820 1.185 ;
        RECT  1.895 0.770 3.340 0.930 ;
        RECT  1.735 0.535 1.895 0.930 ;
        RECT  0.735 0.535 1.735 0.695 ;
        RECT  0.575 0.535 0.735 1.225 ;
        RECT  0.340 0.965 0.575 1.225 ;
        END
        AntennaGateArea 0.2366 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.410 3.375 1.630 ;
        RECT  2.470 1.320 2.850 1.630 ;
        RECT  1.030 1.470 2.470 1.630 ;
        RECT  0.770 1.440 1.030 1.630 ;
        END
        AntennaGateArea 0.2366 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 2.250 2.895 2.410 ;
        RECT  1.235 2.150 1.655 2.410 ;
        END
        AntennaGateArea 0.2366 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.460 1.110 2.200 1.270 ;
        RECT  1.280 0.880 1.460 1.270 ;
        RECT  0.920 0.880 1.280 1.170 ;
        END
        AntennaGateArea 0.2366 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 -0.130 5.330 0.130 ;
        RECT  4.945 -0.130 5.205 0.980 ;
        RECT  4.075 -0.130 4.945 0.130 ;
        RECT  3.815 -0.130 4.075 0.250 ;
        RECT  0.385 -0.130 3.815 0.130 ;
        RECT  0.125 -0.130 0.385 0.755 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 2.740 5.330 3.000 ;
        RECT  4.945 1.860 5.205 3.000 ;
        RECT  4.125 2.740 4.945 3.000 ;
        RECT  3.865 2.570 4.125 3.000 ;
        RECT  3.605 2.740 3.865 3.000 ;
        RECT  3.005 2.570 3.605 3.000 ;
        RECT  2.470 2.740 3.005 3.000 ;
        RECT  1.870 2.620 2.470 3.000 ;
        RECT  1.545 2.740 1.870 3.000 ;
        RECT  0.945 2.620 1.545 3.000 ;
        RECT  0.725 2.740 0.945 3.000 ;
        RECT  0.125 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.275 1.225 4.305 1.485 ;
        RECT  4.115 0.430 4.275 1.970 ;
        RECT  2.085 0.430 4.115 0.590 ;
        RECT  0.535 1.810 4.115 1.970 ;
    END
END AND4X4MTH

MACRO AND4X6MTH
    CLASS CORE ;
    FOREIGN AND4X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.995 0.385 7.255 2.410 ;
        RECT  6.175 1.290 6.995 1.580 ;
        RECT  5.915 0.385 6.175 2.410 ;
        END
        AntennaDiffArea 1.143 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.275 1.135 1.580 ;
        END
        AntennaGateArea 0.286 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.515 1.275 2.170 1.580 ;
        END
        AntennaGateArea 0.286 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.175 1.275 3.725 1.580 ;
        END
        AntennaGateArea 0.286 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.275 4.750 1.580 ;
        END
        AntennaGateArea 0.286 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.710 -0.130 7.380 0.130 ;
        RECT  6.450 -0.130 6.710 1.000 ;
        RECT  5.610 -0.130 6.450 0.130 ;
        RECT  5.350 -0.130 5.610 1.000 ;
        RECT  0.935 -0.130 5.350 0.130 ;
        RECT  0.675 -0.130 0.935 0.640 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.715 2.740 7.380 3.000 ;
        RECT  6.455 1.770 6.715 3.000 ;
        RECT  5.630 2.740 6.455 3.000 ;
        RECT  5.370 1.790 5.630 3.000 ;
        RECT  5.190 2.740 5.370 3.000 ;
        RECT  4.930 2.155 5.190 3.000 ;
        RECT  4.650 2.740 4.930 3.000 ;
        RECT  4.390 2.560 4.650 3.000 ;
        RECT  4.105 2.740 4.390 3.000 ;
        RECT  3.845 2.155 4.105 3.000 ;
        RECT  3.560 2.740 3.845 3.000 ;
        RECT  3.300 2.560 3.560 3.000 ;
        RECT  2.970 2.740 3.300 3.000 ;
        RECT  2.370 2.230 2.970 3.000 ;
        RECT  2.035 2.740 2.370 3.000 ;
        RECT  1.775 2.560 2.035 3.000 ;
        RECT  1.485 2.740 1.775 3.000 ;
        RECT  1.225 2.120 1.485 3.000 ;
        RECT  0.935 2.740 1.225 3.000 ;
        RECT  0.675 2.560 0.935 3.000 ;
        RECT  0.385 2.740 0.675 3.000 ;
        RECT  0.125 1.810 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.165 1.235 5.710 1.495 ;
        RECT  5.005 0.815 5.165 1.930 ;
        RECT  4.075 0.470 5.100 0.630 ;
        RECT  4.325 0.815 5.005 0.975 ;
        RECT  4.645 1.770 5.005 1.930 ;
        RECT  4.385 1.770 4.645 2.030 ;
        RECT  3.555 1.770 4.385 1.930 ;
        RECT  3.815 0.470 4.075 0.975 ;
        RECT  2.775 0.815 3.815 0.975 ;
        RECT  3.295 0.385 3.555 0.630 ;
        RECT  3.295 1.770 3.555 2.030 ;
        RECT  2.005 0.385 3.295 0.545 ;
        RECT  2.035 1.770 3.295 1.930 ;
        RECT  2.265 0.750 2.525 1.015 ;
        RECT  1.485 0.855 2.265 1.015 ;
        RECT  1.775 1.770 2.035 2.030 ;
        RECT  1.745 0.385 2.005 0.675 ;
        RECT  0.935 1.770 1.775 1.930 ;
        RECT  1.225 0.415 1.485 1.015 ;
        RECT  0.385 0.855 1.225 1.015 ;
        RECT  0.675 1.770 0.935 2.030 ;
        RECT  0.125 0.415 0.385 1.015 ;
    END
END AND4X6MTH

MACRO AND4X8MTH
    CLASS CORE ;
    FOREIGN AND4X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.725 1.685 1.985 2.410 ;
        RECT  1.710 0.385 1.780 0.985 ;
        RECT  1.710 1.685 1.725 2.035 ;
        RECT  1.360 0.385 1.710 2.035 ;
        RECT  0.925 1.085 1.360 1.785 ;
        RECT  0.840 1.085 0.925 2.285 ;
        RECT  0.665 0.385 0.840 2.285 ;
        RECT  0.580 0.385 0.665 1.785 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 1.275 3.495 1.560 ;
        END
        AntennaGateArea 0.4251 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.855 1.275 4.895 1.560 ;
        END
        AntennaGateArea 0.4251 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.605 1.280 6.545 1.560 ;
        END
        AntennaGateArea 0.4251 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.055 1.280 7.995 1.580 ;
        END
        AntennaGateArea 0.4251 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 -0.130 8.610 0.130 ;
        RECT  2.060 -0.130 2.320 0.980 ;
        RECT  0.000 -0.130 2.060 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.485 2.740 8.610 3.000 ;
        RECT  8.225 2.130 8.485 3.000 ;
        RECT  7.885 2.740 8.225 3.000 ;
        RECT  7.285 2.570 7.885 3.000 ;
        RECT  6.935 2.740 7.285 3.000 ;
        RECT  6.335 2.570 6.935 3.000 ;
        RECT  5.905 2.740 6.335 3.000 ;
        RECT  5.305 2.570 5.905 3.000 ;
        RECT  4.865 2.740 5.305 3.000 ;
        RECT  4.265 2.570 4.865 3.000 ;
        RECT  3.905 2.740 4.265 3.000 ;
        RECT  3.305 2.570 3.905 3.000 ;
        RECT  2.865 2.740 3.305 3.000 ;
        RECT  2.265 2.570 2.865 3.000 ;
        RECT  1.455 2.740 2.265 3.000 ;
        RECT  1.195 2.255 1.455 3.000 ;
        RECT  0.385 2.740 1.195 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.380 0.740 8.485 1.020 ;
        RECT  8.225 0.740 8.380 1.940 ;
        RECT  8.220 0.860 8.225 1.940 ;
        RECT  7.465 0.860 8.220 1.020 ;
        RECT  2.325 1.780 8.220 1.940 ;
        RECT  7.715 0.455 7.975 0.675 ;
        RECT  6.950 0.455 7.715 0.615 ;
        RECT  7.205 0.815 7.465 1.020 ;
        RECT  6.690 0.455 6.950 0.725 ;
        RECT  5.910 0.455 6.690 0.615 ;
        RECT  6.170 0.815 6.430 1.025 ;
        RECT  5.390 0.865 6.170 1.025 ;
        RECT  5.650 0.455 5.910 0.675 ;
        RECT  5.130 0.750 5.390 1.025 ;
        RECT  4.350 0.865 5.130 1.025 ;
        RECT  4.610 0.450 4.870 0.685 ;
        RECT  3.830 0.450 4.610 0.610 ;
        RECT  4.090 0.815 4.350 1.025 ;
        RECT  3.570 0.450 3.830 0.840 ;
        RECT  2.610 0.580 3.570 0.840 ;
        RECT  2.165 1.235 2.325 1.940 ;
        RECT  1.895 1.235 2.165 1.495 ;
    END
END AND4X8MTH

MACRO AND4XLMTH
    CLASS CORE ;
    FOREIGN AND4XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.765 2.770 2.195 ;
        RECT  2.485 0.765 2.610 1.175 ;
        RECT  2.485 1.935 2.610 2.195 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.720 0.765 1.960 1.395 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.445 1.540 0.760 ;
        END
        AntennaGateArea 0.0533 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.805 1.300 1.130 1.990 ;
        END
        AntennaGateArea 0.0533 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.535 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 -0.130 2.870 0.130 ;
        RECT  1.920 -0.130 2.520 0.515 ;
        RECT  1.610 -0.130 1.920 0.130 ;
        RECT  1.010 -0.130 1.610 0.250 ;
        RECT  0.730 -0.130 1.010 0.130 ;
        RECT  0.130 -0.130 0.730 0.300 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.465 2.740 2.870 3.000 ;
        RECT  1.865 2.620 2.465 3.000 ;
        RECT  1.640 2.740 1.865 3.000 ;
        RECT  1.040 2.620 1.640 3.000 ;
        RECT  0.000 2.740 1.040 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.170 1.495 2.400 1.755 ;
        RECT  1.740 1.595 2.170 1.755 ;
        RECT  1.480 1.595 1.740 2.400 ;
        RECT  1.470 1.595 1.480 1.755 ;
        RECT  0.790 2.240 1.480 2.400 ;
        RECT  1.310 0.940 1.470 1.755 ;
        RECT  0.385 0.940 1.310 1.100 ;
        RECT  0.530 2.215 0.790 2.400 ;
        RECT  0.125 0.765 0.385 1.100 ;
    END
END AND4XLMTH

MACRO ANTENNAMTH
    CLASS CORE ANTENNACELL ;
    FOREIGN ANTENNAMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.820 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.280 0.645 0.540 2.300 ;
        RECT  0.100 1.290 0.280 1.580 ;
        END
        AntennaDiffArea 0.72590 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 -0.130 0.820 0.130 ;
        RECT  0.280 -0.130 0.540 0.300 ;
        RECT  0.000 -0.130 0.280 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.740 0.820 3.000 ;
        RECT  0.280 2.570 0.540 3.000 ;
        RECT  0.000 2.740 0.280 3.000 ;
        END
    END VDD
END ANTENNAMTH

MACRO AO21X1MTH
    CLASS CORE ;
    FOREIGN AO21X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 1.290 2.770 1.580 ;
        RECT  2.485 0.725 2.745 2.230 ;
        RECT  2.225 0.725 2.485 0.985 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.205 1.680 1.580 ;
        END
        AntennaGateArea 0.065 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.625 1.585 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.810 1.205 1.130 1.620 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 -0.130 2.870 0.130 ;
        RECT  1.665 -0.130 1.925 0.590 ;
        RECT  1.300 -0.130 1.665 0.130 ;
        RECT  0.800 -0.130 1.300 0.340 ;
        RECT  0.465 -0.130 0.800 0.130 ;
        RECT  0.205 -0.130 0.465 0.975 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 2.740 2.870 3.000 ;
        RECT  1.945 2.265 2.205 3.000 ;
        RECT  1.615 2.740 1.945 3.000 ;
        RECT  0.675 2.490 1.615 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.025 1.225 2.265 1.485 ;
        RECT  1.865 0.865 2.025 1.950 ;
        RECT  1.355 0.865 1.865 1.025 ;
        RECT  1.575 1.790 1.865 1.950 ;
        RECT  1.095 0.765 1.355 1.025 ;
        RECT  0.125 1.800 1.325 1.960 ;
    END
END AO21X1MTH

MACRO AO21X2MTH
    CLASS CORE ;
    FOREIGN AO21X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 1.290 2.770 1.580 ;
        RECT  2.485 0.395 2.745 2.415 ;
        RECT  2.225 0.395 2.485 0.995 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.205 1.680 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.625 1.585 ;
        END
        AntennaGateArea 0.1144 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.810 1.205 1.130 1.620 ;
        END
        AntennaGateArea 0.1144 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 -0.130 2.870 0.130 ;
        RECT  1.645 -0.130 1.905 0.590 ;
        RECT  1.300 -0.130 1.645 0.130 ;
        RECT  0.800 -0.130 1.300 0.340 ;
        RECT  0.465 -0.130 0.800 0.130 ;
        RECT  0.205 -0.130 0.465 0.975 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 2.740 2.870 3.000 ;
        RECT  1.975 2.185 2.235 3.000 ;
        RECT  1.615 2.740 1.975 3.000 ;
        RECT  0.675 2.490 1.615 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.025 1.225 2.265 1.485 ;
        RECT  1.865 0.865 2.025 1.920 ;
        RECT  1.275 0.865 1.865 1.025 ;
        RECT  1.575 1.760 1.865 1.920 ;
        RECT  1.065 1.800 1.325 2.060 ;
        RECT  1.115 0.765 1.275 1.025 ;
        RECT  0.385 1.800 1.065 1.960 ;
        RECT  0.125 1.800 0.385 2.060 ;
    END
END AO21X2MTH

MACRO AO21X4MTH
    CLASS CORE ;
    FOREIGN AO21X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.090 1.290 3.180 1.580 ;
        RECT  2.910 0.365 3.090 2.415 ;
        RECT  2.715 0.365 2.910 0.965 ;
        RECT  2.785 1.815 2.910 2.415 ;
        END
        AntennaDiffArea 0.636 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.380 1.210 1.990 1.580 ;
        END
        AntennaGateArea 0.1924 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.160 0.585 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.765 1.205 1.185 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 1.025 ;
        RECT  2.290 -0.130 3.305 0.130 ;
        RECT  1.690 -0.130 2.290 0.680 ;
        RECT  0.385 -0.130 1.690 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 2.740 3.690 3.000 ;
        RECT  3.295 1.800 3.555 3.000 ;
        RECT  2.505 2.740 3.295 3.000 ;
        RECT  2.245 2.180 2.505 3.000 ;
        RECT  0.905 2.740 2.245 3.000 ;
        RECT  0.645 2.185 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.530 1.225 2.730 1.485 ;
        RECT  2.370 0.865 2.530 1.935 ;
        RECT  1.245 0.865 2.370 1.025 ;
        RECT  1.955 1.775 2.370 1.935 ;
        RECT  1.695 1.775 1.955 2.440 ;
        RECT  1.165 1.840 1.425 2.440 ;
        RECT  0.985 0.355 1.245 1.025 ;
        RECT  0.385 1.840 1.165 2.000 ;
        RECT  0.125 1.840 0.385 2.440 ;
    END
END AO21X4MTH

MACRO AO21X8MTH
    CLASS CORE ;
    FOREIGN AO21X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.255 0.390 5.515 2.415 ;
        RECT  5.020 0.745 5.255 2.015 ;
        RECT  4.495 0.745 5.020 1.045 ;
        RECT  4.495 1.665 5.020 2.015 ;
        RECT  4.235 0.370 4.495 1.045 ;
        RECT  4.235 1.665 4.495 2.415 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.190 3.135 1.545 ;
        END
        AntennaGateArea 0.3848 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.205 2.145 1.685 ;
        RECT  0.725 1.525 1.885 1.685 ;
        RECT  0.465 1.205 0.725 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.185 1.605 1.345 ;
        RECT  0.920 0.880 1.130 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 -0.130 6.150 0.130 ;
        RECT  5.765 -0.130 6.025 0.955 ;
        RECT  5.005 -0.130 5.765 0.130 ;
        RECT  4.745 -0.130 5.005 0.565 ;
        RECT  3.905 -0.130 4.745 0.130 ;
        RECT  3.305 -0.130 3.905 0.630 ;
        RECT  2.390 -0.130 3.305 0.130 ;
        RECT  2.130 -0.130 2.390 0.630 ;
        RECT  0.585 -0.130 2.130 0.130 ;
        RECT  0.325 -0.130 0.585 0.955 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 2.740 6.150 3.000 ;
        RECT  5.765 1.850 6.025 3.000 ;
        RECT  5.005 2.740 5.765 3.000 ;
        RECT  4.745 2.215 5.005 3.000 ;
        RECT  3.985 2.740 4.745 3.000 ;
        RECT  3.725 1.815 3.985 3.000 ;
        RECT  0.935 2.740 3.725 3.000 ;
        RECT  0.675 2.205 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.545 1.225 4.790 1.485 ;
        RECT  3.385 0.845 3.545 1.885 ;
        RECT  3.215 2.070 3.475 2.465 ;
        RECT  2.965 0.845 3.385 1.005 ;
        RECT  2.955 1.725 3.385 1.885 ;
        RECT  2.435 2.305 3.215 2.465 ;
        RECT  2.705 0.625 2.965 1.005 ;
        RECT  2.695 1.725 2.955 2.080 ;
        RECT  1.480 0.845 2.705 1.005 ;
        RECT  2.175 1.865 2.435 2.465 ;
        RECT  1.485 1.865 2.175 2.025 ;
        RECT  1.225 1.865 1.485 2.465 ;
        RECT  1.320 0.435 1.480 1.005 ;
        RECT  1.185 0.435 1.320 0.695 ;
        RECT  0.385 1.865 1.225 2.025 ;
        RECT  0.125 1.865 0.385 2.465 ;
    END
END AO21X8MTH

MACRO AO21XLMTH
    CLASS CORE ;
    FOREIGN AO21XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 0.635 2.365 2.480 ;
        RECT  2.125 0.635 2.205 0.895 ;
        RECT  2.150 1.700 2.205 2.480 ;
        RECT  2.045 2.220 2.150 2.480 ;
        END
        AntennaDiffArea 0.219 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.120 0.920 1.580 1.380 ;
        END
        AntennaGateArea 0.0533 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 0.880 0.720 1.370 ;
        END
        AntennaGateArea 0.0533 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.770 2.005 1.190 2.360 ;
        END
        AntennaGateArea 0.0533 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 -0.130 2.460 0.130 ;
        RECT  1.530 -0.130 2.130 0.380 ;
        RECT  0.725 -0.130 1.530 0.130 ;
        RECT  0.385 -0.130 0.725 0.355 ;
        RECT  0.125 -0.130 0.385 0.695 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 2.740 2.460 3.000 ;
        RECT  1.505 2.215 1.765 3.000 ;
        RECT  1.315 2.740 1.505 3.000 ;
        RECT  0.375 2.540 1.315 3.000 ;
        RECT  0.000 2.740 0.375 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.965 1.105 2.025 1.365 ;
        RECT  1.945 1.105 1.965 1.905 ;
        RECT  1.785 0.580 1.945 1.905 ;
        RECT  1.015 0.580 1.785 0.740 ;
        RECT  1.705 1.645 1.785 1.905 ;
        RECT  0.385 1.665 1.395 1.825 ;
        RECT  0.125 1.665 0.385 1.945 ;
    END
END AO21XLMTH

MACRO AO22X1MTH
    CLASS CORE ;
    FOREIGN AO22X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 1.700 3.180 2.385 ;
        RECT  2.965 0.455 3.155 2.385 ;
        RECT  2.895 0.455 2.965 0.715 ;
        RECT  2.895 2.125 2.965 2.385 ;
        END
        AntennaDiffArea 0.329 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.970 0.660 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 0.985 1.140 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.140 0.430 2.440 0.965 ;
        END
        AntennaGateArea 0.0598 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 0.960 1.620 1.580 ;
        END
        AntennaGateArea 0.0598 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.525 -0.130 3.280 0.130 ;
        RECT  2.265 -0.130 2.525 0.250 ;
        RECT  0.500 -0.130 2.265 0.130 ;
        RECT  0.240 -0.130 0.500 0.695 ;
        RECT  0.000 -0.130 0.240 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.615 2.740 3.280 3.000 ;
        RECT  2.015 2.480 2.615 3.000 ;
        RECT  1.645 2.740 2.015 3.000 ;
        RECT  0.705 2.480 1.645 3.000 ;
        RECT  0.000 2.740 0.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.620 0.995 2.780 1.305 ;
        RECT  1.960 1.145 2.620 1.305 ;
        RECT  2.510 1.485 2.610 1.645 ;
        RECT  2.350 1.485 2.510 2.195 ;
        RECT  1.520 2.035 2.350 2.195 ;
        RECT  1.960 1.695 2.060 1.855 ;
        RECT  1.800 0.610 1.960 1.855 ;
        RECT  1.390 0.610 1.800 0.770 ;
        RECT  1.760 1.695 1.800 1.855 ;
        RECT  1.360 1.765 1.520 2.195 ;
        RECT  1.130 0.510 1.390 0.770 ;
        RECT  0.125 1.765 1.360 1.925 ;
    END
END AO22X1MTH

MACRO AO22X2MTH
    CLASS CORE ;
    FOREIGN AO22X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 1.290 3.590 2.380 ;
        RECT  3.380 0.425 3.540 2.380 ;
        RECT  3.290 0.425 3.380 1.025 ;
        RECT  3.300 1.780 3.380 2.380 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.100 0.650 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.830 1.090 1.130 1.645 ;
        END
        AntennaGateArea 0.1053 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.160 1.165 2.770 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.085 1.640 1.650 ;
        END
        AntennaGateArea 0.1053 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.860 -0.130 3.690 0.130 ;
        RECT  2.260 -0.130 2.860 0.630 ;
        RECT  1.790 -0.130 2.260 0.130 ;
        RECT  0.850 -0.130 1.790 0.300 ;
        RECT  0.490 -0.130 0.850 0.130 ;
        RECT  0.230 -0.130 0.490 0.910 ;
        RECT  0.000 -0.130 0.230 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 2.740 3.690 3.000 ;
        RECT  2.820 1.835 3.020 3.000 ;
        RECT  2.320 2.740 2.820 3.000 ;
        RECT  1.380 2.570 2.320 3.000 ;
        RECT  0.950 2.740 1.380 3.000 ;
        RECT  0.690 2.240 0.950 3.000 ;
        RECT  0.350 2.530 0.690 3.000 ;
        RECT  0.000 2.740 0.350 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.110 1.235 3.170 1.495 ;
        RECT  2.950 0.825 3.110 1.495 ;
        RECT  1.980 0.825 2.950 0.985 ;
        RECT  2.440 1.875 2.540 2.035 ;
        RECT  2.280 1.875 2.440 2.330 ;
        RECT  1.520 2.170 2.280 2.330 ;
        RECT  1.980 1.830 2.030 1.990 ;
        RECT  1.820 0.745 1.980 1.990 ;
        RECT  1.125 0.745 1.820 0.905 ;
        RECT  1.770 1.830 1.820 1.990 ;
        RECT  1.360 1.830 1.520 2.330 ;
        RECT  0.125 1.830 1.360 1.990 ;
    END
END AO22X2MTH

MACRO AO22X4MTH
    CLASS CORE ;
    FOREIGN AO22X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 1.290 3.590 1.580 ;
        RECT  3.350 0.410 3.530 2.380 ;
        RECT  3.175 0.410 3.350 1.010 ;
        RECT  3.200 1.780 3.350 2.380 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.160 0.615 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.175 1.130 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.175 2.360 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.175 1.770 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.100 0.130 ;
        RECT  3.715 -0.130 3.975 0.995 ;
        RECT  2.815 -0.130 3.715 0.130 ;
        RECT  2.215 -0.130 2.815 0.655 ;
        RECT  0.420 -0.130 2.215 0.130 ;
        RECT  0.160 -0.130 0.420 0.975 ;
        RECT  0.000 -0.130 0.160 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 2.740 4.100 3.000 ;
        RECT  3.710 1.835 3.970 3.000 ;
        RECT  0.935 2.740 3.710 3.000 ;
        RECT  0.675 2.115 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.985 1.240 3.170 1.500 ;
        RECT  2.825 0.835 2.985 1.920 ;
        RECT  1.395 0.835 2.825 0.995 ;
        RECT  1.995 1.760 2.825 1.920 ;
        RECT  2.245 2.110 2.505 2.395 ;
        RECT  1.485 2.235 2.245 2.395 ;
        RECT  1.735 1.760 1.995 2.020 ;
        RECT  1.225 1.760 1.485 2.395 ;
        RECT  1.135 0.395 1.395 0.995 ;
        RECT  0.385 1.760 1.225 1.920 ;
        RECT  0.125 1.760 0.385 2.380 ;
    END
END AO22X4MTH

MACRO AO22X8MTH
    CLASS CORE ;
    FOREIGN AO22X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.075 0.405 6.335 2.415 ;
        RECT  5.840 0.745 6.075 2.120 ;
        RECT  5.315 0.745 5.840 1.045 ;
        RECT  5.355 1.770 5.840 2.120 ;
        RECT  5.095 1.770 5.355 2.415 ;
        RECT  5.055 0.405 5.315 1.045 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 1.245 2.085 1.685 ;
        RECT  0.785 1.525 1.825 1.685 ;
        RECT  0.435 1.135 0.785 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.185 1.590 1.345 ;
        RECT  0.985 0.880 1.540 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.835 1.295 3.995 1.695 ;
        RECT  2.770 1.535 3.835 1.695 ;
        RECT  2.450 1.225 2.770 1.695 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 0.880 3.565 1.355 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 -0.130 6.970 0.130 ;
        RECT  6.585 -0.130 6.845 0.955 ;
        RECT  5.825 -0.130 6.585 0.130 ;
        RECT  5.565 -0.130 5.825 0.565 ;
        RECT  4.705 -0.130 5.565 0.130 ;
        RECT  4.105 -0.130 4.705 0.765 ;
        RECT  2.340 -0.130 4.105 0.130 ;
        RECT  2.080 -0.130 2.340 0.695 ;
        RECT  0.585 -0.130 2.080 0.130 ;
        RECT  0.325 -0.130 0.585 0.920 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 1.815 6.845 3.000 ;
        RECT  4.815 2.740 6.585 3.000 ;
        RECT  4.655 1.735 4.815 3.000 ;
        RECT  4.555 1.735 4.655 1.895 ;
        RECT  0.905 2.740 4.655 3.000 ;
        RECT  0.645 2.230 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.335 1.225 5.570 1.485 ;
        RECT  4.155 2.245 4.415 2.465 ;
        RECT  4.175 0.950 4.335 2.065 ;
        RECT  3.925 0.950 4.175 1.110 ;
        RECT  2.595 1.905 4.175 2.065 ;
        RECT  2.375 2.245 4.155 2.405 ;
        RECT  3.765 0.540 3.925 1.110 ;
        RECT  2.690 0.540 3.765 0.700 ;
        RECT  2.530 0.540 2.690 1.045 ;
        RECT  1.900 0.885 2.530 1.045 ;
        RECT  2.115 1.875 2.375 2.475 ;
        RECT  1.425 1.875 2.115 2.035 ;
        RECT  1.740 0.505 1.900 1.045 ;
        RECT  1.115 0.505 1.740 0.665 ;
        RECT  1.165 1.875 1.425 2.475 ;
        RECT  0.385 1.875 1.165 2.035 ;
        RECT  0.125 1.875 0.385 2.475 ;
    END
END AO22X8MTH

MACRO AO22XLMTH
    CLASS CORE ;
    FOREIGN AO22XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 1.700 3.180 2.385 ;
        RECT  2.965 0.625 3.155 2.385 ;
        RECT  2.895 0.625 2.965 0.885 ;
        RECT  2.895 2.125 2.965 2.385 ;
        END
        AntennaDiffArea 0.234 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.100 0.660 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.000 1.240 1.140 1.585 ;
        RECT  0.840 0.845 1.000 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 0.405 2.110 0.720 ;
        END
        AntennaGateArea 0.0533 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.600 1.240 1.700 1.515 ;
        RECT  1.320 1.240 1.600 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.900 -0.130 3.280 0.130 ;
        RECT  2.560 -0.130 2.900 0.305 ;
        RECT  2.300 -0.130 2.560 0.880 ;
        RECT  1.300 -0.130 2.300 0.130 ;
        RECT  0.700 -0.130 1.300 0.305 ;
        RECT  0.500 -0.130 0.700 0.130 ;
        RECT  0.240 -0.130 0.500 0.915 ;
        RECT  0.000 -0.130 0.240 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.615 2.740 3.280 3.000 ;
        RECT  2.015 2.375 2.615 3.000 ;
        RECT  1.645 2.740 2.015 3.000 ;
        RECT  0.705 2.480 1.645 3.000 ;
        RECT  0.000 2.740 0.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.040 1.185 2.765 1.445 ;
        RECT  2.380 1.625 2.610 1.785 ;
        RECT  2.220 1.625 2.380 2.195 ;
        RECT  1.600 2.035 2.220 2.195 ;
        RECT  1.880 0.900 2.040 1.855 ;
        RECT  1.340 0.900 1.880 1.060 ;
        RECT  1.780 1.695 1.880 1.855 ;
        RECT  1.440 1.765 1.600 2.195 ;
        RECT  0.125 1.765 1.440 1.925 ;
        RECT  1.180 0.655 1.340 1.060 ;
    END
END AO22XLMTH

MACRO AO2B2BX1MTH
    CLASS CORE ;
    FOREIGN AO2B2BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 0.665 4.820 2.430 ;
        RECT  4.535 0.665 4.610 0.925 ;
        RECT  4.535 2.170 4.610 2.430 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.215 0.720 2.045 ;
        END
        AntennaGateArea 0.0546 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.660 0.985 1.960 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.875 1.565 4.410 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.140 0.960 2.440 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 -0.130 4.920 0.130 ;
        RECT  3.995 -0.130 4.255 0.250 ;
        RECT  3.175 -0.130 3.995 0.130 ;
        RECT  2.915 -0.130 3.175 0.250 ;
        RECT  1.305 -0.130 2.915 0.130 ;
        RECT  0.705 -0.130 1.305 0.695 ;
        RECT  0.000 -0.130 0.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 2.740 4.920 3.000 ;
        RECT  3.995 2.530 4.255 3.000 ;
        RECT  1.280 2.740 3.995 3.000 ;
        RECT  1.280 2.225 1.635 2.485 ;
        RECT  1.020 2.225 1.280 3.000 ;
        RECT  0.695 2.225 1.020 2.485 ;
        RECT  0.000 2.740 1.020 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.355 1.095 4.405 1.355 ;
        RECT  4.195 0.430 4.355 1.355 ;
        RECT  2.785 0.430 4.195 0.590 ;
        RECT  3.535 1.425 3.695 2.485 ;
        RECT  3.125 0.775 3.685 0.935 ;
        RECT  3.125 1.425 3.535 1.585 ;
        RECT  3.185 1.765 3.355 1.925 ;
        RECT  3.025 1.765 3.185 2.265 ;
        RECT  2.965 0.775 3.125 1.585 ;
        RECT  2.340 2.105 3.025 2.265 ;
        RECT  2.625 0.430 2.785 1.925 ;
        RECT  2.210 0.430 2.625 0.590 ;
        RECT  2.525 1.765 2.625 1.925 ;
        RECT  2.180 1.765 2.340 2.265 ;
        RECT  1.950 0.430 2.210 0.775 ;
        RECT  0.900 1.765 2.180 1.925 ;
        RECT  1.315 0.875 1.475 1.585 ;
        RECT  0.335 0.875 1.315 1.035 ;
        RECT  0.330 2.155 0.360 2.415 ;
        RECT  0.330 0.515 0.335 1.035 ;
        RECT  0.170 0.515 0.330 2.415 ;
    END
END AO2B2BX1MTH

MACRO AO2B2BX2MTH
    CLASS CORE ;
    FOREIGN AO2B2BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 0.380 4.820 2.405 ;
        RECT  4.535 0.380 4.610 0.980 ;
        RECT  4.535 1.805 4.610 2.405 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.215 0.720 2.045 ;
        END
        AntennaGateArea 0.0546 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.660 0.985 1.960 1.585 ;
        END
        AntennaGateArea 0.1053 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.155 4.000 1.835 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.140 0.960 2.435 1.585 ;
        END
        AntennaGateArea 0.1053 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 -0.130 4.920 0.130 ;
        RECT  3.995 -0.130 4.255 0.250 ;
        RECT  3.175 -0.130 3.995 0.130 ;
        RECT  2.915 -0.130 3.175 0.250 ;
        RECT  1.305 -0.130 2.915 0.130 ;
        RECT  0.705 -0.130 1.305 0.695 ;
        RECT  0.000 -0.130 0.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 2.740 4.920 3.000 ;
        RECT  4.025 2.015 4.285 3.000 ;
        RECT  1.635 2.740 4.025 3.000 ;
        RECT  0.695 2.485 1.635 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.355 1.135 4.405 1.395 ;
        RECT  4.195 0.430 4.355 1.395 ;
        RECT  2.775 0.430 4.195 0.590 ;
        RECT  3.610 2.015 3.715 2.175 ;
        RECT  3.115 0.815 3.685 0.975 ;
        RECT  3.450 1.425 3.610 2.175 ;
        RECT  3.115 1.425 3.450 1.585 ;
        RECT  2.995 1.765 3.155 2.265 ;
        RECT  2.955 0.815 3.115 1.585 ;
        RECT  2.185 2.105 2.995 2.265 ;
        RECT  2.615 0.430 2.775 1.925 ;
        RECT  2.210 0.430 2.615 0.590 ;
        RECT  2.435 1.765 2.615 1.925 ;
        RECT  1.950 0.430 2.210 0.775 ;
        RECT  2.025 1.765 2.185 2.265 ;
        RECT  0.900 1.765 2.025 1.925 ;
        RECT  1.315 0.875 1.475 1.585 ;
        RECT  0.335 0.875 1.315 1.035 ;
        RECT  0.330 2.155 0.360 2.415 ;
        RECT  0.330 0.515 0.335 1.035 ;
        RECT  0.170 0.515 0.330 2.415 ;
    END
END AO2B2BX2MTH

MACRO AO2B2BX4MTH
    CLASS CORE ;
    FOREIGN AO2B2BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.985 0.355 5.175 2.300 ;
        RECT  4.845 0.355 4.985 0.955 ;
        RECT  4.845 1.700 4.985 2.300 ;
        RECT  4.610 1.700 4.845 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.215 0.925 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.070 1.085 2.370 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.100 1.575 4.425 1.990 ;
        END
        AntennaGateArea 0.0897 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 1.085 2.770 1.685 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 0.955 ;
        RECT  4.565 -0.130 5.355 0.130 ;
        RECT  4.305 -0.130 4.565 0.250 ;
        RECT  3.485 -0.130 4.305 0.130 ;
        RECT  3.225 -0.130 3.485 0.250 ;
        RECT  1.435 -0.130 3.225 0.130 ;
        RECT  0.835 -0.130 1.435 0.695 ;
        RECT  0.000 -0.130 0.835 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 1.700 5.615 3.000 ;
        RECT  4.595 2.740 5.355 3.000 ;
        RECT  4.335 2.170 4.595 3.000 ;
        RECT  2.035 2.740 4.335 3.000 ;
        RECT  1.775 2.220 2.035 3.000 ;
        RECT  0.925 2.740 1.775 3.000 ;
        RECT  0.665 1.805 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.665 1.135 4.805 1.395 ;
        RECT  4.505 0.430 4.665 1.395 ;
        RECT  3.110 0.430 4.505 0.590 ;
        RECT  3.920 2.170 4.085 2.330 ;
        RECT  3.450 0.815 4.030 0.975 ;
        RECT  3.760 1.425 3.920 2.330 ;
        RECT  3.450 1.425 3.760 1.585 ;
        RECT  3.365 1.765 3.525 2.365 ;
        RECT  3.290 0.815 3.450 1.585 ;
        RECT  2.555 2.205 3.365 2.365 ;
        RECT  2.950 0.430 3.110 2.025 ;
        RECT  2.520 0.430 2.950 0.590 ;
        RECT  2.805 1.865 2.950 2.025 ;
        RECT  2.395 1.870 2.555 2.365 ;
        RECT  2.260 0.405 2.520 0.905 ;
        RECT  1.520 1.870 2.395 2.030 ;
        RECT  1.445 1.155 1.785 1.415 ;
        RECT  1.260 1.760 1.520 2.360 ;
        RECT  1.285 0.875 1.445 1.415 ;
        RECT  0.415 0.875 1.285 1.035 ;
        RECT  0.315 0.765 0.415 1.035 ;
        RECT  0.315 1.760 0.415 1.920 ;
        RECT  0.155 0.765 0.315 1.920 ;
    END
END AO2B2BX4MTH

MACRO AO2B2BXLMTH
    CLASS CORE ;
    FOREIGN AO2B2BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 0.725 4.820 2.330 ;
        RECT  4.585 0.725 4.610 0.985 ;
        RECT  4.535 2.170 4.610 2.330 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN B1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.215 0.720 2.045 ;
        END
        AntennaGateArea 0.0546 ;
    END B1N
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.660 0.985 1.960 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.875 1.575 4.410 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.140 0.960 2.440 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 -0.130 4.920 0.130 ;
        RECT  3.995 -0.130 4.255 0.250 ;
        RECT  3.175 -0.130 3.995 0.130 ;
        RECT  2.915 -0.130 3.175 0.250 ;
        RECT  1.305 -0.130 2.915 0.130 ;
        RECT  0.705 -0.130 1.305 0.695 ;
        RECT  0.000 -0.130 0.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 2.740 4.920 3.000 ;
        RECT  3.995 2.580 4.255 3.000 ;
        RECT  1.280 2.740 3.995 3.000 ;
        RECT  1.280 2.225 1.635 2.485 ;
        RECT  1.020 2.225 1.280 3.000 ;
        RECT  0.695 2.225 1.020 2.485 ;
        RECT  0.000 2.740 1.020 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.355 1.095 4.405 1.355 ;
        RECT  4.195 0.430 4.355 1.355 ;
        RECT  2.785 0.430 4.195 0.590 ;
        RECT  3.535 1.425 3.695 2.485 ;
        RECT  3.125 0.775 3.685 0.935 ;
        RECT  3.125 1.425 3.535 1.585 ;
        RECT  3.185 1.765 3.355 1.925 ;
        RECT  3.025 1.765 3.185 2.265 ;
        RECT  2.965 0.775 3.125 1.585 ;
        RECT  2.340 2.105 3.025 2.265 ;
        RECT  2.625 0.430 2.785 1.925 ;
        RECT  2.210 0.430 2.625 0.590 ;
        RECT  2.525 1.765 2.625 1.925 ;
        RECT  2.180 1.765 2.340 2.265 ;
        RECT  2.000 0.430 2.210 0.775 ;
        RECT  0.900 1.765 2.180 1.925 ;
        RECT  1.950 0.515 2.000 0.775 ;
        RECT  1.315 0.875 1.475 1.585 ;
        RECT  0.335 0.875 1.315 1.035 ;
        RECT  0.330 2.155 0.360 2.415 ;
        RECT  0.330 0.515 0.335 1.035 ;
        RECT  0.170 0.515 0.330 2.415 ;
    END
END AO2B2BXLMTH

MACRO AO2B2X1MTH
    CLASS CORE ;
    FOREIGN AO2B2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.665 4.000 2.430 ;
        RECT  3.715 0.665 3.790 0.925 ;
        RECT  3.715 2.170 3.790 2.430 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.970 0.660 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 0.985 1.140 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.055 1.565 3.590 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 0.960 1.620 1.585 ;
        END
        AntennaGateArea 0.0598 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 -0.130 4.100 0.130 ;
        RECT  3.175 -0.130 3.435 0.250 ;
        RECT  2.355 -0.130 3.175 0.130 ;
        RECT  2.095 -0.130 2.355 0.250 ;
        RECT  0.495 -0.130 2.095 0.130 ;
        RECT  0.235 -0.130 0.495 0.695 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  3.175 2.530 3.435 3.000 ;
        RECT  0.965 2.740 3.175 3.000 ;
        RECT  0.705 2.195 0.965 3.000 ;
        RECT  0.000 2.740 0.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.535 1.095 3.585 1.355 ;
        RECT  3.375 0.430 3.535 1.355 ;
        RECT  1.965 0.430 3.375 0.590 ;
        RECT  2.715 1.425 2.875 2.485 ;
        RECT  2.305 0.775 2.865 0.935 ;
        RECT  2.305 1.425 2.715 1.585 ;
        RECT  2.365 1.765 2.535 1.925 ;
        RECT  2.205 1.765 2.365 2.265 ;
        RECT  2.145 0.775 2.305 1.585 ;
        RECT  1.520 2.105 2.205 2.265 ;
        RECT  1.805 0.430 1.965 1.925 ;
        RECT  1.390 0.430 1.805 0.590 ;
        RECT  1.705 1.765 1.805 1.925 ;
        RECT  1.360 1.765 1.520 2.265 ;
        RECT  1.130 0.430 1.390 0.775 ;
        RECT  0.125 1.765 1.360 1.925 ;
    END
END AO2B2X1MTH

MACRO AO2B2X2MTH
    CLASS CORE ;
    FOREIGN AO2B2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.425 4.000 2.340 ;
        RECT  3.765 0.425 3.790 1.025 ;
        RECT  3.715 1.740 3.790 2.340 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.970 0.660 1.585 ;
        END
        AntennaGateArea 0.1053 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 0.985 1.140 1.585 ;
        END
        AntennaGateArea 0.1053 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.185 3.245 1.815 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 0.985 1.615 1.585 ;
        END
        AntennaGateArea 0.1053 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 -0.130 4.100 0.130 ;
        RECT  3.175 -0.130 3.435 0.250 ;
        RECT  2.355 -0.130 3.175 0.130 ;
        RECT  2.095 -0.130 2.355 0.250 ;
        RECT  0.495 -0.130 2.095 0.130 ;
        RECT  0.235 -0.130 0.495 0.790 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 2.740 4.100 3.000 ;
        RECT  3.205 1.995 3.465 3.000 ;
        RECT  0.935 2.740 3.205 3.000 ;
        RECT  0.675 2.385 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.425 0.430 3.585 1.395 ;
        RECT  1.955 0.430 3.425 0.590 ;
        RECT  2.295 0.815 2.865 0.975 ;
        RECT  2.790 1.995 2.845 2.255 ;
        RECT  2.630 1.425 2.790 2.255 ;
        RECT  2.295 1.425 2.630 1.585 ;
        RECT  2.175 1.765 2.335 2.265 ;
        RECT  2.135 0.815 2.295 1.585 ;
        RECT  1.365 2.105 2.175 2.265 ;
        RECT  1.795 0.430 1.955 1.925 ;
        RECT  1.425 0.430 1.795 0.590 ;
        RECT  1.615 1.765 1.795 1.925 ;
        RECT  1.165 0.430 1.425 0.805 ;
        RECT  1.205 1.765 1.365 2.265 ;
        RECT  0.130 1.765 1.205 1.925 ;
    END
END AO2B2X2MTH

MACRO AO2B2X4MTH
    CLASS CORE ;
    FOREIGN AO2B2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.710 0.380 3.900 2.385 ;
        RECT  3.665 0.380 3.710 0.980 ;
        RECT  3.615 1.700 3.710 2.385 ;
        RECT  3.380 1.700 3.615 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.970 0.660 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 1.110 1.140 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.185 3.020 1.580 ;
        END
        AntennaGateArea 0.0884 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 1.110 1.615 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  4.125 -0.130 4.385 0.980 ;
        RECT  3.335 -0.130 4.125 0.130 ;
        RECT  3.075 -0.130 3.335 0.250 ;
        RECT  2.355 -0.130 3.075 0.130 ;
        RECT  2.095 -0.130 2.355 0.250 ;
        RECT  0.495 -0.130 2.095 0.130 ;
        RECT  0.235 -0.130 0.495 0.790 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.785 4.385 3.000 ;
        RECT  3.335 2.740 4.125 3.000 ;
        RECT  3.075 2.325 3.335 3.000 ;
        RECT  0.905 2.740 3.075 3.000 ;
        RECT  0.645 2.105 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.485 1.135 3.530 1.395 ;
        RECT  3.325 0.430 3.485 1.395 ;
        RECT  1.955 0.430 3.325 0.590 ;
        RECT  2.295 1.760 2.895 1.920 ;
        RECT  2.295 0.815 2.865 0.975 ;
        RECT  2.235 2.205 2.395 2.515 ;
        RECT  2.135 0.815 2.295 1.920 ;
        RECT  1.425 2.205 2.235 2.365 ;
        RECT  1.795 0.430 1.955 1.925 ;
        RECT  1.390 0.430 1.795 0.590 ;
        RECT  1.675 1.765 1.795 1.925 ;
        RECT  1.165 1.765 1.425 2.365 ;
        RECT  1.130 0.430 1.390 0.930 ;
        RECT  0.390 1.765 1.165 1.925 ;
        RECT  0.130 1.765 0.390 2.365 ;
    END
END AO2B2X4MTH

MACRO AO2B2XLMTH
    CLASS CORE ;
    FOREIGN AO2B2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.620 4.000 2.330 ;
        RECT  3.765 0.620 3.790 0.880 ;
        RECT  3.715 2.170 3.790 2.330 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.970 0.660 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 0.985 1.140 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.055 1.475 3.590 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 0.960 1.620 1.585 ;
        END
        AntennaGateArea 0.0533 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 -0.130 4.100 0.130 ;
        RECT  3.175 -0.130 3.435 0.250 ;
        RECT  2.355 -0.130 3.175 0.130 ;
        RECT  2.095 -0.130 2.355 0.250 ;
        RECT  0.495 -0.130 2.095 0.130 ;
        RECT  0.235 -0.130 0.495 0.775 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  3.175 2.580 3.435 3.000 ;
        RECT  0.965 2.740 3.175 3.000 ;
        RECT  0.705 2.195 0.965 3.000 ;
        RECT  0.000 2.740 0.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.535 0.995 3.585 1.255 ;
        RECT  3.375 0.430 3.535 1.255 ;
        RECT  1.965 0.430 3.375 0.590 ;
        RECT  2.715 1.425 2.875 2.485 ;
        RECT  2.305 0.780 2.865 0.940 ;
        RECT  2.305 1.425 2.715 1.585 ;
        RECT  2.365 1.765 2.535 1.925 ;
        RECT  2.205 1.765 2.365 2.265 ;
        RECT  2.145 0.780 2.305 1.585 ;
        RECT  1.520 2.105 2.205 2.265 ;
        RECT  1.805 0.430 1.965 1.925 ;
        RECT  1.390 0.430 1.805 0.590 ;
        RECT  1.705 1.765 1.805 1.925 ;
        RECT  1.360 1.765 1.520 2.265 ;
        RECT  1.130 0.430 1.390 0.770 ;
        RECT  0.125 1.765 1.360 1.925 ;
    END
END AO2B2XLMTH

MACRO AOI211X1MTH
    CLASS CORE ;
    FOREIGN AOI211X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.540 2.360 2.125 ;
        RECT  1.810 0.540 2.200 0.700 ;
        RECT  2.150 1.700 2.200 2.125 ;
        RECT  1.980 1.865 2.150 2.125 ;
        RECT  1.550 0.540 1.810 0.915 ;
        RECT  0.125 0.540 1.550 0.700 ;
        END
        AntennaDiffArea 0.471 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 1.095 1.540 1.675 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.095 2.020 1.500 ;
        RECT  1.720 1.095 1.950 1.685 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 0.880 1.050 1.540 ;
        RECT  0.510 0.880 0.785 1.170 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.350 0.565 1.690 ;
        RECT  0.100 1.290 0.310 1.690 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  2.075 -0.130 2.335 0.300 ;
        RECT  1.600 -0.130 2.075 0.130 ;
        RECT  1.000 -0.130 1.600 0.300 ;
        RECT  0.000 -0.130 1.000 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 2.740 2.460 3.000 ;
        RECT  1.325 2.555 2.265 3.000 ;
        RECT  1.100 2.740 1.325 3.000 ;
        RECT  0.160 2.555 1.100 3.000 ;
        RECT  0.000 2.740 0.160 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.150 1.875 1.410 2.135 ;
        RECT  0.385 1.875 1.150 2.035 ;
        RECT  0.125 1.875 0.385 2.135 ;
    END
END AOI211X1MTH

MACRO AOI211X2MTH
    CLASS CORE ;
    FOREIGN AOI211X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 0.755 2.365 2.500 ;
        RECT  1.815 0.755 2.205 0.915 ;
        RECT  2.150 1.700 2.205 2.500 ;
        RECT  1.985 1.900 2.150 2.500 ;
        RECT  1.555 0.415 1.815 0.915 ;
        RECT  0.385 0.540 1.555 0.700 ;
        RECT  0.125 0.440 0.385 0.700 ;
        END
        AntennaDiffArea 0.811 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.230 1.095 1.545 1.660 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.095 2.025 1.500 ;
        RECT  1.725 1.095 1.950 1.685 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 0.880 1.050 1.540 ;
        RECT  0.510 0.880 0.785 1.170 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.350 0.565 1.690 ;
        RECT  0.100 1.290 0.310 1.690 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  2.075 -0.130 2.335 0.575 ;
        RECT  1.265 -0.130 2.075 0.130 ;
        RECT  1.005 -0.130 1.265 0.360 ;
        RECT  0.000 -0.130 1.005 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 2.740 2.460 3.000 ;
        RECT  0.645 2.220 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.165 1.875 1.425 2.475 ;
        RECT  0.385 1.875 1.165 2.035 ;
        RECT  0.125 1.875 0.385 2.475 ;
    END
END AOI211X2MTH

MACRO AOI211X4MTH
    CLASS CORE ;
    FOREIGN AOI211X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.850 0.540 4.010 2.125 ;
        RECT  0.955 0.540 3.850 0.800 ;
        RECT  3.790 1.540 3.850 2.125 ;
        RECT  2.895 1.865 3.790 2.125 ;
        END
        AntennaDiffArea 1.074 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.510 0.980 3.670 1.345 ;
        RECT  2.495 0.980 3.510 1.140 ;
        RECT  2.150 0.980 2.495 1.660 ;
        END
        AntennaGateArea 0.3796 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.710 1.330 3.225 1.670 ;
        END
        AntennaGateArea 0.3796 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 0.990 1.965 1.595 ;
        RECT  0.555 0.990 1.700 1.150 ;
        RECT  0.295 0.990 0.555 1.455 ;
        END
        AntennaGateArea 0.3926 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.330 1.395 1.540 ;
        END
        AntennaGateArea 0.3926 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.035 -0.130 4.100 0.130 ;
        RECT  2.775 -0.130 3.035 0.360 ;
        RECT  0.385 -0.130 2.775 0.130 ;
        RECT  0.125 -0.130 0.385 0.800 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 2.740 4.100 3.000 ;
        RECT  1.565 2.220 1.825 3.000 ;
        RECT  0.000 2.740 1.565 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.335 2.305 3.975 2.465 ;
        RECT  2.075 1.875 2.335 2.465 ;
        RECT  1.315 1.875 2.075 2.035 ;
        RECT  1.055 1.875 1.315 2.475 ;
        RECT  0.385 1.875 1.055 2.035 ;
        RECT  0.125 1.875 0.385 2.475 ;
    END
END AOI211X4MTH

MACRO AOI211XLMTH
    CLASS CORE ;
    FOREIGN AOI211XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.540 2.370 2.060 ;
        RECT  1.800 0.540 2.210 0.700 ;
        RECT  2.150 1.700 2.210 2.060 ;
        RECT  1.990 1.830 2.150 2.060 ;
        RECT  1.540 0.540 1.800 0.915 ;
        RECT  0.125 0.540 1.540 0.700 ;
        END
        AntennaDiffArea 0.36 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.205 1.095 1.550 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.095 2.030 1.500 ;
        RECT  1.730 1.095 1.950 1.650 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 0.880 1.025 1.540 ;
        RECT  0.510 0.880 0.785 1.170 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.350 0.595 1.580 ;
        RECT  0.100 1.075 0.310 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  1.735 -0.130 2.335 0.300 ;
        RECT  1.525 -0.130 1.735 0.130 ;
        RECT  0.685 -0.130 1.525 0.300 ;
        RECT  0.000 -0.130 0.685 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 2.740 2.460 3.000 ;
        RECT  1.550 2.570 2.150 3.000 ;
        RECT  1.275 2.740 1.550 3.000 ;
        RECT  0.335 2.335 1.275 3.000 ;
        RECT  0.000 2.740 0.335 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.125 1.770 1.420 1.930 ;
    END
END AOI211XLMTH

MACRO AOI21BX1MTH
    CLASS CORE ;
    FOREIGN AOI21BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.730 2.770 2.115 ;
        RECT  2.485 0.730 2.610 0.990 ;
        RECT  2.485 1.700 2.610 2.115 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 2.125 2.060 2.360 ;
        END
        AntennaGateArea 0.078 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.765 2.080 1.275 2.360 ;
        END
        AntennaGateArea 0.0572 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.975 0.460 1.580 ;
        END
        AntennaGateArea 0.0572 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 -0.130 2.870 0.130 ;
        RECT  1.605 -0.130 2.205 0.475 ;
        RECT  0.385 -0.130 1.605 0.130 ;
        RECT  0.125 -0.130 0.385 0.565 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 2.740 2.870 3.000 ;
        RECT  1.265 2.540 2.205 3.000 ;
        RECT  1.065 2.740 1.265 3.000 ;
        RECT  0.125 2.540 1.065 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.305 1.225 2.430 1.485 ;
        RECT  2.145 0.865 2.305 1.845 ;
        RECT  1.495 0.865 2.145 1.025 ;
        RECT  1.795 1.685 2.145 1.845 ;
        RECT  1.535 1.685 1.795 1.945 ;
        RECT  0.985 1.225 1.625 1.485 ;
        RECT  1.235 0.765 1.495 1.025 ;
        RECT  0.825 0.355 0.985 1.895 ;
        RECT  0.725 0.355 0.825 0.515 ;
        RECT  0.565 1.735 0.825 1.895 ;
    END
END AOI21BX1MTH

MACRO AOI21BX2MTH
    CLASS CORE ;
    FOREIGN AOI21BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.390 2.770 2.370 ;
        RECT  2.485 0.390 2.610 0.990 ;
        RECT  2.485 1.700 2.610 2.370 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 2.125 2.175 2.360 ;
        END
        AntennaGateArea 0.0962 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 2.080 1.275 2.360 ;
        END
        AntennaGateArea 0.0572 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.970 0.445 1.580 ;
        END
        AntennaGateArea 0.0572 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 -0.130 2.870 0.130 ;
        RECT  1.605 -0.130 2.205 0.405 ;
        RECT  0.385 -0.130 1.605 0.130 ;
        RECT  0.125 -0.130 0.385 0.565 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 2.740 2.870 3.000 ;
        RECT  1.265 2.540 2.205 3.000 ;
        RECT  1.065 2.740 1.265 3.000 ;
        RECT  0.125 2.540 1.065 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.305 1.225 2.405 1.485 ;
        RECT  2.145 0.865 2.305 1.845 ;
        RECT  1.495 0.865 2.145 1.025 ;
        RECT  1.795 1.685 2.145 1.845 ;
        RECT  1.535 1.685 1.795 1.945 ;
        RECT  0.985 1.225 1.625 1.485 ;
        RECT  1.235 0.765 1.495 1.025 ;
        RECT  0.825 0.355 0.985 1.895 ;
        RECT  0.725 0.355 0.825 0.515 ;
        RECT  0.565 1.735 0.825 1.895 ;
    END
END AOI21BX2MTH

MACRO AOI21BX4MTH
    CLASS CORE ;
    FOREIGN AOI21BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.370 0.825 3.590 1.955 ;
        RECT  3.025 0.825 3.370 1.045 ;
        RECT  3.025 1.735 3.370 1.955 ;
        RECT  2.765 0.390 3.025 1.045 ;
        RECT  2.765 1.735 3.025 2.435 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.205 2.225 1.580 ;
        END
        AntennaGateArea 0.1885 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.115 1.205 1.580 ;
        END
        AntennaGateArea 0.0884 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.875 0.355 1.695 ;
        END
        AntennaGateArea 0.0884 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.630 ;
        RECT  2.485 -0.130 3.305 0.130 ;
        RECT  2.225 -0.130 2.485 0.630 ;
        RECT  1.065 -0.130 2.225 0.130 ;
        RECT  0.125 -0.130 1.065 0.435 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 2.740 3.690 3.000 ;
        RECT  3.305 2.165 3.565 3.000 ;
        RECT  2.485 2.740 3.305 3.000 ;
        RECT  2.225 2.100 2.485 3.000 ;
        RECT  1.370 2.740 2.225 3.000 ;
        RECT  1.110 2.140 1.370 3.000 ;
        RECT  0.725 2.740 1.110 3.000 ;
        RECT  0.125 2.280 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.565 1.245 3.145 1.505 ;
        RECT  2.405 0.835 2.565 1.920 ;
        RECT  1.625 0.835 2.405 0.995 ;
        RECT  1.885 1.760 2.405 1.920 ;
        RECT  1.725 1.760 1.885 2.360 ;
        RECT  1.365 0.395 1.625 0.995 ;
        RECT  1.385 1.235 1.545 1.935 ;
        RECT  0.695 1.775 1.385 1.935 ;
        RECT  0.695 0.775 1.115 0.935 ;
        RECT  0.535 0.775 0.695 1.935 ;
    END
END AOI21BX4MTH

MACRO AOI21BX8MTH
    CLASS CORE ;
    FOREIGN AOI21BX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.435 0.390 4.695 2.435 ;
        RECT  4.200 0.745 4.435 2.120 ;
        RECT  3.675 0.745 4.200 1.085 ;
        RECT  3.765 1.780 4.200 2.120 ;
        RECT  3.505 1.780 3.765 2.435 ;
        RECT  3.415 0.390 3.675 1.085 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.160 2.875 1.695 ;
        RECT  1.515 1.535 2.560 1.695 ;
        RECT  1.355 1.195 1.515 1.695 ;
        END
        AntennaGateArea 0.377 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.195 0.355 1.910 ;
        END
        AntennaGateArea 0.1781 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.165 1.170 1.660 ;
        END
        AntennaGateArea 0.1781 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 -0.130 5.330 0.130 ;
        RECT  4.945 -0.130 5.205 0.990 ;
        RECT  4.185 -0.130 4.945 0.130 ;
        RECT  3.925 -0.130 4.185 0.565 ;
        RECT  3.120 -0.130 3.925 0.130 ;
        RECT  2.860 -0.130 3.120 0.640 ;
        RECT  1.315 -0.130 2.860 0.130 ;
        RECT  1.020 -0.130 1.315 0.640 ;
        RECT  0.000 -0.130 1.020 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 2.740 5.330 3.000 ;
        RECT  4.945 1.835 5.205 3.000 ;
        RECT  3.255 2.740 4.945 3.000 ;
        RECT  2.995 2.265 3.255 3.000 ;
        RECT  1.305 2.740 2.995 3.000 ;
        RECT  1.045 1.875 1.305 3.000 ;
        RECT  0.000 2.740 1.045 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.230 1.265 3.935 1.525 ;
        RECT  3.070 0.820 3.230 2.035 ;
        RECT  2.290 0.820 3.070 0.980 ;
        RECT  2.745 1.875 3.070 2.035 ;
        RECT  2.485 1.875 2.745 2.475 ;
        RECT  1.815 1.875 2.485 2.035 ;
        RECT  1.945 1.165 2.360 1.355 ;
        RECT  2.130 0.380 2.290 0.980 ;
        RECT  1.955 0.380 2.130 0.640 ;
        RECT  1.785 0.825 1.945 1.355 ;
        RECT  1.555 1.875 1.815 2.475 ;
        RECT  0.695 0.825 1.785 0.985 ;
        RECT  0.695 1.825 0.765 2.425 ;
        RECT  0.535 0.825 0.695 2.425 ;
        RECT  0.385 0.825 0.535 0.985 ;
        RECT  0.125 0.385 0.385 0.985 ;
    END
END AOI21BX8MTH

MACRO AOI21BXLMTH
    CLASS CORE ;
    FOREIGN AOI21BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.335 2.770 1.990 ;
        RECT  2.485 0.335 2.610 0.595 ;
        RECT  2.485 1.700 2.610 1.990 ;
        END
        AntennaDiffArea 0.339 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 2.125 2.060 2.360 ;
        END
        AntennaGateArea 0.078 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.765 2.080 1.275 2.360 ;
        END
        AntennaGateArea 0.0572 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.975 0.460 1.580 ;
        END
        AntennaGateArea 0.0572 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 -0.130 2.870 0.130 ;
        RECT  1.605 -0.130 2.205 0.475 ;
        RECT  0.385 -0.130 1.605 0.130 ;
        RECT  0.125 -0.130 0.385 0.545 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 2.740 2.870 3.000 ;
        RECT  1.265 2.540 2.205 3.000 ;
        RECT  1.065 2.740 1.265 3.000 ;
        RECT  0.125 2.540 1.065 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.305 1.225 2.405 1.485 ;
        RECT  2.145 0.865 2.305 1.845 ;
        RECT  1.495 0.865 2.145 1.025 ;
        RECT  1.795 1.685 2.145 1.845 ;
        RECT  1.535 1.685 1.795 1.945 ;
        RECT  0.985 1.225 1.625 1.485 ;
        RECT  1.235 0.765 1.495 1.025 ;
        RECT  0.825 0.355 0.985 1.895 ;
        RECT  0.725 0.355 0.825 0.515 ;
        RECT  0.565 1.735 0.825 1.895 ;
    END
END AOI21BXLMTH

MACRO AOI21X1MTH
    CLASS CORE ;
    FOREIGN AOI21X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.290 1.950 2.085 ;
        RECT  1.740 0.770 1.900 2.085 ;
        RECT  0.985 0.770 1.740 0.930 ;
        RECT  1.665 1.825 1.740 2.085 ;
        END
        AntennaDiffArea 0.347 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.110 1.560 1.645 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.545 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 1.110 1.130 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 -0.130 2.050 0.130 ;
        RECT  1.525 -0.130 1.785 0.590 ;
        RECT  1.270 -0.130 1.525 0.130 ;
        RECT  0.670 -0.130 1.270 0.380 ;
        RECT  0.385 -0.130 0.670 0.130 ;
        RECT  0.125 -0.130 0.385 1.000 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.865 2.740 2.050 3.000 ;
        RECT  1.265 2.620 1.865 3.000 ;
        RECT  1.085 2.740 1.265 3.000 ;
        RECT  0.145 2.620 1.085 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.155 1.880 1.415 2.140 ;
        RECT  0.425 1.880 1.155 2.040 ;
        RECT  0.165 1.880 0.425 2.140 ;
    END
END AOI21X1MTH

MACRO AOI21X2MTH
    CLASS CORE ;
    FOREIGN AOI21X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.290 1.950 2.450 ;
        RECT  1.740 0.795 1.900 2.450 ;
        RECT  1.245 0.795 1.740 0.955 ;
        RECT  1.665 1.850 1.740 2.450 ;
        RECT  0.985 0.355 1.245 0.955 ;
        END
        AntennaDiffArea 0.566 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.135 1.560 1.670 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.210 0.595 1.655 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.775 1.135 1.130 1.660 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.795 -0.130 2.050 0.130 ;
        RECT  1.535 -0.130 1.795 0.615 ;
        RECT  0.385 -0.130 1.535 0.130 ;
        RECT  0.125 -0.130 0.385 1.005 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 2.740 2.050 3.000 ;
        RECT  0.645 2.190 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.155 1.850 1.415 2.450 ;
        RECT  0.385 1.850 1.155 2.010 ;
        RECT  0.125 1.850 0.385 2.450 ;
    END
END AOI21X2MTH

MACRO AOI21X3MTH
    CLASS CORE ;
    FOREIGN AOI21X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.170 1.290 3.295 1.580 ;
        RECT  3.010 0.865 3.170 2.155 ;
        RECT  2.970 0.620 3.010 2.155 ;
        RECT  2.750 0.620 2.970 1.065 ;
        RECT  2.795 1.825 2.970 2.155 ;
        RECT  1.995 0.865 2.750 1.065 ;
        RECT  1.795 0.500 1.995 1.065 ;
        RECT  1.190 0.500 1.795 0.700 ;
        END
        AntennaDiffArea 0.71 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.245 2.790 1.580 ;
        END
        AntennaGateArea 0.312 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.250 2.075 1.685 ;
        RECT  0.730 1.525 1.915 1.685 ;
        RECT  0.465 1.200 0.730 1.685 ;
        END
        AntennaGateArea 0.312 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.000 0.880 1.600 1.345 ;
        END
        AntennaGateArea 0.312 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.675 ;
        RECT  2.445 -0.130 3.305 0.130 ;
        RECT  2.185 -0.130 2.445 0.675 ;
        RECT  0.560 -0.130 2.185 0.130 ;
        RECT  0.300 -0.130 0.560 0.945 ;
        RECT  0.000 -0.130 0.300 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 2.740 3.690 3.000 ;
        RECT  1.750 2.205 2.010 3.000 ;
        RECT  0.925 2.740 1.750 3.000 ;
        RECT  0.665 2.205 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.355 1.810 3.515 2.520 ;
        RECT  2.545 2.360 3.355 2.520 ;
        RECT  2.285 1.865 2.545 2.520 ;
        RECT  1.465 1.865 2.285 2.025 ;
        RECT  1.205 1.865 1.465 2.365 ;
        RECT  0.385 1.865 1.205 2.025 ;
        RECT  0.125 1.865 0.385 2.365 ;
    END
END AOI21X3MTH

MACRO AOI21X4MTH
    CLASS CORE ;
    FOREIGN AOI21X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.170 1.290 3.270 1.580 ;
        RECT  2.985 0.865 3.170 2.155 ;
        RECT  2.970 0.405 2.985 2.155 ;
        RECT  2.725 0.405 2.970 1.065 ;
        RECT  2.795 1.795 2.970 2.155 ;
        RECT  1.980 0.865 2.725 1.065 ;
        RECT  1.780 0.465 1.980 1.065 ;
        RECT  1.190 0.465 1.780 0.665 ;
        END
        AntennaDiffArea 0.908 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.255 2.790 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.250 2.075 1.685 ;
        RECT  0.730 1.525 1.915 1.685 ;
        RECT  0.465 1.205 0.730 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.000 0.880 1.600 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.675 ;
        RECT  2.420 -0.130 3.305 0.130 ;
        RECT  2.160 -0.130 2.420 0.675 ;
        RECT  0.600 -0.130 2.160 0.130 ;
        RECT  0.340 -0.130 0.600 1.025 ;
        RECT  0.000 -0.130 0.340 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 2.740 3.690 3.000 ;
        RECT  1.750 2.205 2.010 3.000 ;
        RECT  0.925 2.740 1.750 3.000 ;
        RECT  0.665 2.205 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.355 1.865 3.515 2.520 ;
        RECT  2.545 2.360 3.355 2.520 ;
        RECT  2.285 1.865 2.545 2.520 ;
        RECT  1.465 1.865 2.285 2.025 ;
        RECT  1.205 1.865 1.465 2.465 ;
        RECT  0.385 1.865 1.205 2.025 ;
        RECT  0.125 1.865 0.385 2.465 ;
    END
END AOI21X4MTH

MACRO AOI21X6MTH
    CLASS CORE ;
    FOREIGN AOI21X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.700 0.405 4.795 1.005 ;
        RECT  4.700 1.760 4.795 2.360 ;
        RECT  4.535 0.405 4.700 2.360 ;
        RECT  4.200 0.800 4.535 2.035 ;
        RECT  3.775 0.800 4.200 1.070 ;
        RECT  3.510 1.765 4.200 2.035 ;
        RECT  3.515 0.405 3.775 1.070 ;
        RECT  3.505 0.540 3.515 1.070 ;
        RECT  0.230 0.540 3.505 0.810 ;
        END
        AntennaDiffArea 1.718 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.325 1.255 3.895 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.725 1.365 2.985 1.685 ;
        RECT  1.605 1.525 2.725 1.685 ;
        RECT  0.980 1.330 1.605 1.685 ;
        END
        AntennaGateArea 0.6162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.805 0.990 2.405 1.345 ;
        RECT  0.720 0.990 1.805 1.150 ;
        RECT  0.375 0.990 0.720 1.585 ;
        END
        AntennaGateArea 0.6162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 -0.130 4.920 0.130 ;
        RECT  4.025 -0.130 4.285 0.615 ;
        RECT  3.220 -0.130 4.025 0.130 ;
        RECT  2.960 -0.130 3.220 0.355 ;
        RECT  1.375 -0.130 2.960 0.130 ;
        RECT  1.115 -0.130 1.375 0.350 ;
        RECT  0.000 -0.130 1.115 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 2.740 4.920 3.000 ;
        RECT  1.565 2.255 1.825 3.000 ;
        RECT  0.000 2.740 1.565 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.265 2.305 4.285 2.465 ;
        RECT  3.005 1.865 3.265 2.465 ;
        RECT  2.335 1.865 3.005 2.025 ;
        RECT  2.075 1.865 2.335 2.465 ;
        RECT  1.315 1.865 2.075 2.025 ;
        RECT  1.055 1.865 1.315 2.465 ;
        RECT  0.385 1.865 1.055 2.025 ;
        RECT  0.125 1.865 0.385 2.465 ;
    END
END AOI21X6MTH

MACRO AOI21X8MTH
    CLASS CORE ;
    FOREIGN AOI21X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 1.165 6.355 1.665 ;
        RECT  5.665 0.405 5.925 2.035 ;
        RECT  5.550 0.800 5.665 2.035 ;
        RECT  4.905 0.800 5.550 1.070 ;
        RECT  4.620 1.765 5.550 2.035 ;
        RECT  4.645 0.405 4.905 1.070 ;
        RECT  4.635 0.540 4.645 1.070 ;
        RECT  1.310 0.540 4.635 0.810 ;
        END
        AntennaDiffArea 1.878 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.465 1.255 5.365 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.835 1.365 4.095 1.685 ;
        RECT  2.630 1.525 3.835 1.685 ;
        RECT  1.985 1.330 2.630 1.685 ;
        RECT  0.725 1.525 1.985 1.685 ;
        RECT  0.465 1.245 0.725 1.685 ;
        END
        AntennaGateArea 0.8216 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.015 0.990 3.615 1.345 ;
        RECT  1.595 0.990 3.015 1.150 ;
        RECT  1.130 0.990 1.595 1.345 ;
        RECT  0.920 0.875 1.130 1.345 ;
        END
        AntennaGateArea 0.8216 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.955 ;
        RECT  5.415 -0.130 6.175 0.130 ;
        RECT  5.155 -0.130 5.415 0.615 ;
        RECT  4.335 -0.130 5.155 0.130 ;
        RECT  4.075 -0.130 4.335 0.355 ;
        RECT  2.460 -0.130 4.075 0.130 ;
        RECT  2.200 -0.130 2.460 0.350 ;
        RECT  0.585 -0.130 2.200 0.130 ;
        RECT  0.325 -0.130 0.585 0.975 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.915 2.740 6.560 3.000 ;
        RECT  2.655 2.205 2.915 3.000 ;
        RECT  0.905 2.740 2.655 3.000 ;
        RECT  0.645 2.205 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.175 1.865 6.435 2.465 ;
        RECT  4.395 2.305 6.175 2.465 ;
        RECT  4.135 1.865 4.395 2.465 ;
        RECT  3.435 1.865 4.135 2.025 ;
        RECT  3.175 1.865 3.435 2.465 ;
        RECT  2.395 1.865 3.175 2.025 ;
        RECT  2.135 1.865 2.395 2.465 ;
        RECT  1.425 1.865 2.135 2.025 ;
        RECT  1.165 1.865 1.425 2.490 ;
        RECT  0.385 1.865 1.165 2.025 ;
        RECT  0.125 1.865 0.385 2.465 ;
    END
END AOI21X8MTH

MACRO AOI21XLMTH
    CLASS CORE ;
    FOREIGN AOI21XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.770 1.950 1.985 ;
        RECT  1.015 0.770 1.740 0.930 ;
        RECT  1.665 1.825 1.740 1.985 ;
        END
        AntennaDiffArea 0.25 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.110 1.560 1.645 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.545 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.730 1.110 1.130 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 -0.130 2.050 0.130 ;
        RECT  1.585 -0.130 1.845 0.590 ;
        RECT  1.270 -0.130 1.585 0.130 ;
        RECT  0.670 -0.130 1.270 0.380 ;
        RECT  0.385 -0.130 0.670 0.130 ;
        RECT  0.125 -0.130 0.385 1.000 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 2.740 2.050 3.000 ;
        RECT  1.200 2.570 1.800 3.000 ;
        RECT  0.965 2.740 1.200 3.000 ;
        RECT  0.365 2.330 0.965 3.000 ;
        RECT  0.000 2.740 0.365 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.165 1.825 1.415 1.985 ;
    END
END AOI21XLMTH

MACRO AOI221X1MTH
    CLASS CORE ;
    FOREIGN AOI221X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.020 0.525 3.180 2.425 ;
        RECT  0.125 0.525 3.020 0.685 ;
        RECT  2.895 1.700 3.020 2.425 ;
        END
        AntennaDiffArea 0.479 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 0.865 2.815 1.325 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.330 1.045 1.605 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 0.865 0.565 1.150 ;
        RECT  0.100 0.865 0.310 1.200 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 0.880 1.525 1.260 ;
        RECT  0.880 0.880 1.265 1.150 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 0.865 2.205 1.325 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 -0.130 3.280 0.130 ;
        RECT  2.485 -0.130 3.085 0.345 ;
        RECT  1.295 -0.130 2.485 0.130 ;
        RECT  1.035 -0.130 1.295 0.345 ;
        RECT  0.000 -0.130 1.035 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.135 2.740 3.280 3.000 ;
        RECT  0.195 2.555 1.135 3.000 ;
        RECT  0.000 2.740 0.195 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.670 2.265 2.610 2.525 ;
        RECT  2.045 1.510 2.305 1.945 ;
        RECT  1.345 1.785 2.045 1.945 ;
        RECT  0.125 1.785 1.345 2.045 ;
    END
END AOI221X1MTH

MACRO AOI221X2MTH
    CLASS CORE ;
    FOREIGN AOI221X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.385 0.815 3.590 2.405 ;
        RECT  3.380 0.375 3.385 2.405 ;
        RECT  3.125 0.375 3.380 0.975 ;
        RECT  3.255 1.805 3.380 2.405 ;
        RECT  1.870 0.815 3.125 0.975 ;
        RECT  1.270 0.375 1.870 0.975 ;
        END
        AntennaDiffArea 1.201 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.810 1.165 3.180 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.160 0.725 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.170 1.395 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.160 2.625 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.595 1.160 1.965 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.835 -0.130 3.690 0.130 ;
        RECT  2.575 -0.130 2.835 0.630 ;
        RECT  0.555 -0.130 2.575 0.130 ;
        RECT  0.295 -0.130 0.555 0.980 ;
        RECT  0.000 -0.130 0.295 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 2.740 3.690 3.000 ;
        RECT  1.195 2.105 1.455 3.000 ;
        RECT  0.385 2.740 1.195 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.745 1.805 3.005 2.560 ;
        RECT  1.975 2.400 2.745 2.560 ;
        RECT  2.225 1.765 2.485 2.220 ;
        RECT  0.905 1.765 2.225 1.925 ;
        RECT  1.715 2.135 1.975 2.560 ;
        RECT  0.645 1.765 0.905 2.400 ;
    END
END AOI221X2MTH

MACRO AOI221X4MTH
    CLASS CORE ;
    FOREIGN AOI221X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.515 0.820 5.640 2.035 ;
        RECT  5.455 0.820 5.515 2.125 ;
        RECT  5.430 0.360 5.455 2.125 ;
        RECT  5.195 0.360 5.430 1.000 ;
        RECT  5.255 1.760 5.430 2.125 ;
        RECT  3.905 0.560 5.195 0.740 ;
        RECT  3.645 0.480 3.905 0.740 ;
        RECT  1.635 0.560 3.645 0.740 ;
        RECT  1.035 0.480 1.635 0.740 ;
        END
        AntennaDiffArea 1.454 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.805 1.205 5.250 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.020 0.990 2.310 1.345 ;
        RECT  0.660 0.990 2.020 1.150 ;
        RECT  0.100 0.990 0.660 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.845 1.330 1.635 1.615 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.365 0.920 4.625 1.465 ;
        RECT  3.265 0.920 4.365 1.080 ;
        RECT  2.930 0.920 3.265 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 1.260 4.125 1.670 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.995 -0.130 6.150 0.130 ;
        RECT  5.735 -0.130 5.995 0.640 ;
        RECT  4.890 -0.130 5.735 0.130 ;
        RECT  4.630 -0.130 4.890 0.380 ;
        RECT  2.935 -0.130 4.630 0.130 ;
        RECT  2.335 -0.130 2.935 0.380 ;
        RECT  0.385 -0.130 2.335 0.130 ;
        RECT  0.125 -0.130 0.385 0.800 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.525 2.740 6.150 3.000 ;
        RECT  2.265 2.300 2.525 3.000 ;
        RECT  1.455 2.740 2.265 3.000 ;
        RECT  1.195 2.200 1.455 3.000 ;
        RECT  0.385 2.740 1.195 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.765 2.205 6.025 2.465 ;
        RECT  5.005 2.305 5.765 2.465 ;
        RECT  4.745 1.795 5.005 2.465 ;
        RECT  2.925 2.305 4.745 2.465 ;
        RECT  4.225 1.865 4.485 2.125 ;
        RECT  3.445 1.865 4.225 2.025 ;
        RECT  3.345 1.865 3.445 2.125 ;
        RECT  3.185 1.525 3.345 2.125 ;
        RECT  1.975 1.525 3.185 1.685 ;
        RECT  2.765 1.865 2.925 2.465 ;
        RECT  2.665 1.865 2.765 2.025 ;
        RECT  1.815 1.525 1.975 2.395 ;
        RECT  1.715 1.795 1.815 2.395 ;
        RECT  0.935 1.795 1.715 1.955 ;
        RECT  0.675 1.795 0.935 2.395 ;
    END
END AOI221X4MTH

MACRO AOI221XLMTH
    CLASS CORE ;
    FOREIGN AOI221XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.620 0.525 2.780 2.425 ;
        RECT  0.125 0.525 2.620 0.685 ;
        RECT  2.485 1.700 2.620 2.425 ;
        END
        AntennaDiffArea 0.377 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.865 2.440 1.465 ;
        END
        AntennaGateArea 0.0702 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.330 1.065 1.605 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 0.865 0.585 1.150 ;
        RECT  0.100 0.865 0.310 1.235 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 0.880 1.530 1.150 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 0.865 1.970 1.465 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 2.870 0.130 ;
        RECT  2.485 -0.130 2.745 0.345 ;
        RECT  1.640 -0.130 2.485 0.130 ;
        RECT  0.700 -0.130 1.640 0.345 ;
        RECT  0.000 -0.130 0.700 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 2.740 2.870 3.000 ;
        RECT  1.055 2.385 1.315 3.000 ;
        RECT  0.795 2.740 1.055 3.000 ;
        RECT  0.195 2.385 0.795 3.000 ;
        RECT  0.000 2.740 0.195 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.045 1.645 2.305 1.955 ;
        RECT  1.635 2.165 2.235 2.425 ;
        RECT  0.125 1.795 2.045 1.955 ;
    END
END AOI221XLMTH

MACRO AOI222X1MTH
    CLASS CORE ;
    FOREIGN AOI222X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.465 3.590 1.935 ;
        RECT  0.125 0.465 3.380 0.625 ;
        RECT  3.055 1.775 3.380 1.935 ;
        RECT  2.795 1.775 3.055 2.220 ;
        END
        AntennaDiffArea 0.632 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 1.330 1.050 1.600 ;
        END
        AntennaGateArea 0.1274 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 0.805 0.575 1.095 ;
        RECT  0.100 0.805 0.310 1.170 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 0.805 1.475 1.130 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 0.865 2.195 1.310 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.810 3.200 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.455 0.835 2.770 1.450 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 -0.130 3.690 0.130 ;
        RECT  3.145 -0.130 3.405 0.250 ;
        RECT  1.295 -0.130 3.145 0.130 ;
        RECT  1.035 -0.130 1.295 0.250 ;
        RECT  0.000 -0.130 1.035 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.075 2.740 3.690 3.000 ;
        RECT  0.135 2.570 1.075 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.305 2.160 3.565 2.560 ;
        RECT  2.355 2.400 3.305 2.560 ;
        RECT  1.755 2.265 2.355 2.560 ;
        RECT  1.995 1.490 2.255 1.945 ;
        RECT  1.315 1.785 1.995 1.945 ;
        RECT  1.055 1.785 1.315 2.045 ;
        RECT  0.385 1.785 1.055 1.945 ;
        RECT  0.125 1.785 0.385 2.045 ;
    END
END AOI222X1MTH

MACRO AOI222X2MTH
    CLASS CORE ;
    FOREIGN AOI222X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.715 0.395 3.975 1.020 ;
        RECT  3.590 0.820 3.715 1.020 ;
        RECT  3.545 0.820 3.590 1.170 ;
        RECT  3.375 0.820 3.545 2.145 ;
        RECT  1.870 0.820 3.375 1.020 ;
        RECT  3.205 1.885 3.375 2.145 ;
        RECT  1.270 0.370 1.870 1.020 ;
        END
        AntennaDiffArea 1.189 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.675 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 1.200 1.285 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 1.200 2.575 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 1.200 1.950 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.215 3.195 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.725 1.290 4.000 1.760 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.115 -0.130 4.100 0.130 ;
        RECT  2.515 -0.130 3.115 0.600 ;
        RECT  0.555 -0.130 2.515 0.130 ;
        RECT  0.295 -0.130 0.555 0.980 ;
        RECT  0.000 -0.130 0.295 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 4.100 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.765 1.940 3.925 2.560 ;
        RECT  2.955 2.400 3.765 2.560 ;
        RECT  2.695 1.805 2.955 2.560 ;
        RECT  1.905 2.400 2.695 2.560 ;
        RECT  2.175 1.765 2.435 2.220 ;
        RECT  0.905 1.765 2.175 1.925 ;
        RECT  1.645 2.135 1.905 2.560 ;
        RECT  0.645 1.765 0.905 2.400 ;
    END
END AOI222X2MTH

MACRO AOI222X4MTH
    CLASS CORE ;
    FOREIGN AOI222X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.630 0.395 6.870 2.085 ;
        RECT  6.385 0.395 6.630 0.995 ;
        RECT  6.335 1.865 6.630 2.085 ;
        RECT  4.700 0.560 6.385 0.740 ;
        RECT  6.075 1.865 6.335 2.220 ;
        RECT  5.315 1.865 6.075 2.085 ;
        RECT  5.055 1.865 5.315 2.215 ;
        RECT  4.440 0.355 4.700 0.955 ;
        RECT  2.685 0.560 4.440 0.740 ;
        RECT  2.085 0.370 2.685 0.970 ;
        RECT  0.410 0.560 2.085 0.740 ;
        RECT  0.150 0.355 0.410 0.955 ;
        END
        AntennaDiffArea 2.298 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 0.920 1.505 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.755 1.200 2.060 1.685 ;
        RECT  0.595 1.525 1.755 1.685 ;
        RECT  0.100 1.200 0.595 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.305 0.920 3.920 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.125 1.210 4.430 1.685 ;
        RECT  3.055 1.525 4.125 1.685 ;
        RECT  2.485 1.200 3.055 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.325 0.920 5.925 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.175 1.215 6.450 1.685 ;
        RECT  4.985 1.525 6.175 1.685 ;
        RECT  4.610 1.215 4.985 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.755 -0.130 6.970 0.130 ;
        RECT  5.495 -0.130 5.755 0.380 ;
        RECT  3.745 -0.130 5.495 0.130 ;
        RECT  3.485 -0.130 3.745 0.380 ;
        RECT  1.315 -0.130 3.485 0.130 ;
        RECT  1.055 -0.130 1.315 0.380 ;
        RECT  0.000 -0.130 1.055 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 2.740 6.970 3.000 ;
        RECT  1.065 2.255 1.325 3.000 ;
        RECT  0.000 2.740 1.065 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.585 2.265 6.845 2.560 ;
        RECT  5.825 2.400 6.585 2.560 ;
        RECT  5.565 2.265 5.825 2.560 ;
        RECT  4.805 2.400 5.565 2.560 ;
        RECT  4.545 1.865 4.805 2.560 ;
        RECT  3.785 2.400 4.545 2.560 ;
        RECT  4.035 1.865 4.295 2.125 ;
        RECT  3.275 1.865 4.035 2.025 ;
        RECT  3.525 2.255 3.785 2.560 ;
        RECT  2.765 2.400 3.525 2.560 ;
        RECT  3.015 1.865 3.275 2.125 ;
        RECT  1.845 1.865 3.015 2.025 ;
        RECT  2.505 2.215 2.765 2.560 ;
        RECT  1.585 1.865 1.845 2.465 ;
        RECT  0.805 1.865 1.585 2.025 ;
        RECT  0.545 1.865 0.805 2.465 ;
    END
END AOI222X4MTH

MACRO AOI222XLMTH
    CLASS CORE ;
    FOREIGN AOI222XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.430 3.590 1.920 ;
        RECT  0.125 0.430 3.380 0.610 ;
        RECT  3.055 1.760 3.380 1.920 ;
        RECT  2.795 1.760 3.055 2.220 ;
        END
        AntennaDiffArea 0.421 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.330 1.215 1.540 ;
        END
        AntennaGateArea 0.0702 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 0.795 0.565 1.095 ;
        RECT  0.100 0.795 0.310 1.170 ;
        END
        AntennaGateArea 0.0702 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 0.790 1.560 1.130 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.865 2.195 1.310 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.800 3.200 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.435 0.790 2.790 1.320 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 -0.130 3.690 0.130 ;
        RECT  3.145 -0.130 3.405 0.250 ;
        RECT  1.350 -0.130 3.145 0.130 ;
        RECT  1.090 -0.130 1.350 0.250 ;
        RECT  0.000 -0.130 1.090 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.570 2.740 3.690 3.000 ;
        RECT  1.310 2.570 1.570 3.000 ;
        RECT  1.070 2.740 1.310 3.000 ;
        RECT  0.725 2.060 1.070 3.000 ;
        RECT  0.130 2.570 0.725 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.305 2.100 3.565 2.560 ;
        RECT  2.530 2.400 3.305 2.560 ;
        RECT  1.930 2.070 2.530 2.560 ;
        RECT  2.255 1.505 2.515 1.880 ;
        RECT  1.555 1.720 2.255 1.880 ;
        RECT  1.295 1.720 1.555 2.005 ;
        RECT  0.385 1.720 1.295 1.880 ;
        RECT  0.125 1.720 0.385 2.005 ;
    END
END AOI222XLMTH

MACRO AOI22X1MTH
    CLASS CORE ;
    FOREIGN AOI22X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 0.520 2.360 1.930 ;
        RECT  1.120 0.520 2.180 0.700 ;
        RECT  2.150 1.290 2.180 1.930 ;
        RECT  1.795 1.770 2.150 1.930 ;
        RECT  1.535 1.770 1.795 2.010 ;
        END
        AntennaDiffArea 0.49 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.315 1.365 0.595 1.645 ;
        RECT  0.100 1.205 0.315 1.645 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.775 0.880 1.025 1.250 ;
        RECT  0.510 0.880 0.775 1.170 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 0.880 1.985 1.145 ;
        RECT  1.720 0.880 1.950 1.540 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.205 0.880 1.540 1.575 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.245 -0.130 2.460 0.130 ;
        RECT  1.985 -0.130 2.245 0.335 ;
        RECT  0.385 -0.130 1.985 0.130 ;
        RECT  0.125 -0.130 0.385 0.680 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 2.740 2.460 3.000 ;
        RECT  0.225 2.550 0.825 3.000 ;
        RECT  0.000 2.740 0.225 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.075 2.125 2.335 2.365 ;
        RECT  1.405 2.205 2.075 2.365 ;
        RECT  1.305 2.205 1.405 2.555 ;
        RECT  1.145 1.825 1.305 2.555 ;
        RECT  0.385 1.825 1.145 1.985 ;
        RECT  0.125 1.825 0.385 2.085 ;
    END
END AOI22X1MTH

MACRO AOI22X2MTH
    CLASS CORE ;
    FOREIGN AOI22X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.730 1.290 2.770 1.580 ;
        RECT  2.550 0.770 2.730 2.020 ;
        RECT  1.470 0.770 2.550 0.950 ;
        RECT  1.815 1.780 2.550 2.020 ;
        RECT  1.210 0.405 1.470 0.950 ;
        END
        AntennaDiffArea 0.738 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.145 0.650 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.830 1.135 1.150 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.130 2.370 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.135 1.735 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 -0.130 2.870 0.130 ;
        RECT  2.165 -0.130 2.425 0.590 ;
        RECT  0.510 -0.130 2.165 0.130 ;
        RECT  0.250 -0.130 0.510 0.945 ;
        RECT  0.000 -0.130 0.250 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.995 2.740 2.870 3.000 ;
        RECT  0.735 2.100 0.995 3.000 ;
        RECT  0.000 2.740 0.735 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.325 2.200 2.585 2.460 ;
        RECT  1.565 2.200 2.325 2.360 ;
        RECT  1.305 1.760 1.565 2.360 ;
        RECT  0.420 1.760 1.305 1.920 ;
        RECT  0.160 1.760 0.420 2.360 ;
    END
END AOI22X2MTH

MACRO AOI22X4MTH
    CLASS CORE ;
    FOREIGN AOI22X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.575 0.630 4.820 2.030 ;
        RECT  4.560 0.630 4.575 0.955 ;
        RECT  2.970 1.850 4.575 2.030 ;
        RECT  4.350 0.345 4.560 0.955 ;
        RECT  4.300 0.345 4.350 0.810 ;
        RECT  2.620 0.630 4.300 0.810 ;
        RECT  2.360 0.405 2.620 0.925 ;
        RECT  0.555 0.745 2.360 0.925 ;
        RECT  0.295 0.405 0.555 0.925 ;
        END
        AntennaDiffArea 1.532 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.225 1.885 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.260 1.225 2.330 1.485 ;
        RECT  2.100 1.225 2.260 1.880 ;
        RECT  0.720 1.720 2.100 1.880 ;
        RECT  0.465 1.225 0.720 1.880 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 1.330 3.800 1.560 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.240 4.390 1.500 ;
        RECT  4.000 0.990 4.160 1.500 ;
        RECT  2.960 0.990 4.000 1.150 ;
        RECT  2.800 0.990 2.960 1.580 ;
        RECT  2.555 1.240 2.800 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.635 -0.130 4.920 0.130 ;
        RECT  3.375 -0.130 3.635 0.450 ;
        RECT  1.720 -0.130 3.375 0.130 ;
        RECT  1.120 -0.130 1.720 0.565 ;
        RECT  0.000 -0.130 1.120 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 2.740 4.920 3.000 ;
        RECT  1.905 2.400 2.165 3.000 ;
        RECT  0.985 2.740 1.905 3.000 ;
        RECT  0.725 2.400 0.985 3.000 ;
        RECT  0.000 2.740 0.725 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.720 2.220 4.760 2.380 ;
        RECT  2.460 1.780 2.720 2.380 ;
        RECT  1.555 2.060 2.460 2.220 ;
        RECT  1.295 2.060 1.555 2.320 ;
        RECT  0.385 2.060 1.295 2.220 ;
        RECT  0.125 2.060 0.385 2.320 ;
    END
END AOI22X4MTH

MACRO AOI22XLMTH
    CLASS CORE ;
    FOREIGN AOI22XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.670 2.360 2.010 ;
        RECT  1.290 0.670 2.200 0.890 ;
        RECT  2.150 1.700 2.200 2.010 ;
        RECT  1.655 1.780 2.150 2.010 ;
        RECT  1.130 0.670 1.290 0.950 ;
        END
        AntennaDiffArea 0.276 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.315 1.365 0.595 1.580 ;
        RECT  0.100 1.205 0.315 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.940 1.165 1.030 1.425 ;
        RECT  0.780 0.880 0.940 1.425 ;
        RECT  0.510 0.880 0.780 1.170 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.070 2.020 1.480 ;
        RECT  1.720 1.070 1.950 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.140 1.540 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.280 -0.130 2.460 0.130 ;
        RECT  2.020 -0.130 2.280 0.490 ;
        RECT  1.655 -0.130 2.020 0.130 ;
        RECT  0.715 -0.130 1.655 0.340 ;
        RECT  0.385 -0.130 0.715 0.130 ;
        RECT  0.125 -0.130 0.385 0.680 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.890 2.740 2.460 3.000 ;
        RECT  0.290 2.295 0.890 3.000 ;
        RECT  0.000 2.740 0.290 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.470 2.295 2.265 2.555 ;
        RECT  1.310 1.760 1.470 2.555 ;
        RECT  0.125 1.760 1.310 1.920 ;
    END
END AOI22XLMTH

MACRO AOI2B1X1MTH
    CLASS CORE ;
    FOREIGN AOI2B1X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.770 2.370 2.090 ;
        RECT  1.780 0.770 2.210 0.930 ;
        RECT  2.150 1.700 2.210 2.090 ;
        RECT  2.075 1.875 2.150 2.090 ;
        RECT  1.500 0.565 1.780 0.930 ;
        END
        AntennaDiffArea 0.355 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.115 2.030 1.485 ;
        RECT  1.730 1.115 1.950 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.430 1.010 0.730 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.110 1.550 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 -0.130 2.460 0.130 ;
        RECT  2.070 -0.130 2.330 0.590 ;
        RECT  0.905 -0.130 2.070 0.130 ;
        RECT  0.645 -0.130 0.905 0.300 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.095 2.740 2.460 3.000 ;
        RECT  1.495 2.555 2.095 3.000 ;
        RECT  1.295 2.740 1.495 3.000 ;
        RECT  0.695 2.555 1.295 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.565 1.760 1.825 2.020 ;
        RECT  0.585 1.760 1.565 1.920 ;
        RECT  0.910 0.595 1.070 1.360 ;
        RECT  0.250 0.595 0.910 0.755 ;
        RECT  0.250 2.345 0.385 2.505 ;
        RECT  0.090 0.595 0.250 2.505 ;
    END
END AOI2B1X1MTH

MACRO AOI2B1X2MTH
    CLASS CORE ;
    FOREIGN AOI2B1X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.770 2.770 2.365 ;
        RECT  1.835 0.770 2.560 0.980 ;
        RECT  2.485 1.765 2.560 2.365 ;
        RECT  1.575 0.380 1.835 0.980 ;
        END
        AntennaDiffArea 0.566 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 1.200 2.360 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.155 0.495 1.625 ;
        END
        AntennaGateArea 0.0871 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.200 1.735 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.715 -0.130 2.870 0.130 ;
        RECT  2.115 -0.130 2.715 0.590 ;
        RECT  0.955 -0.130 2.115 0.130 ;
        RECT  0.695 -0.130 0.955 0.590 ;
        RECT  0.355 -0.130 0.695 0.310 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.835 2.740 2.870 3.000 ;
        RECT  1.575 2.265 1.835 3.000 ;
        RECT  0.785 2.740 1.575 3.000 ;
        RECT  0.185 2.315 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.325 1.760 2.235 1.920 ;
        RECT  1.065 1.760 1.325 2.390 ;
        RECT  0.845 1.240 1.105 1.505 ;
        RECT  0.685 0.815 0.845 1.965 ;
        RECT  0.125 0.815 0.685 0.975 ;
        RECT  0.125 1.805 0.685 1.965 ;
    END
END AOI2B1X2MTH

MACRO AOI2B1X4MTH
    CLASS CORE ;
    FOREIGN AOI2B1X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 0.865 4.060 1.580 ;
        RECT  3.825 0.865 3.990 2.155 ;
        RECT  3.790 0.405 3.825 2.155 ;
        RECT  3.565 0.405 3.790 1.065 ;
        RECT  3.610 1.795 3.790 2.155 ;
        RECT  2.810 0.865 3.565 1.065 ;
        RECT  2.610 0.465 2.810 1.065 ;
        RECT  2.005 0.465 2.610 0.665 ;
        END
        AntennaDiffArea 0.912 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.150 1.255 3.605 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.330 1.240 1.005 1.555 ;
        END
        AntennaGateArea 0.1755 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.815 0.880 2.415 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 -0.130 4.510 0.130 ;
        RECT  4.120 -0.130 4.380 0.675 ;
        RECT  3.260 -0.130 4.120 0.130 ;
        RECT  3.000 -0.130 3.260 0.675 ;
        RECT  1.330 -0.130 3.000 0.130 ;
        RECT  0.730 -0.130 1.330 0.720 ;
        RECT  0.000 -0.130 0.730 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 2.740 4.510 3.000 ;
        RECT  2.565 2.205 2.825 3.000 ;
        RECT  0.385 2.740 2.565 3.000 ;
        RECT  0.125 1.830 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.170 1.865 4.390 2.520 ;
        RECT  3.360 2.360 4.170 2.520 ;
        RECT  3.100 1.865 3.360 2.520 ;
        RECT  2.290 1.865 3.100 2.025 ;
        RECT  2.730 1.250 2.890 1.685 ;
        RECT  1.595 1.525 2.730 1.685 ;
        RECT  2.030 1.865 2.290 2.515 ;
        RECT  1.035 2.255 2.030 2.515 ;
        RECT  1.335 0.900 1.595 1.915 ;
        RECT  0.385 0.900 1.335 1.060 ;
        RECT  0.895 1.755 1.335 1.915 ;
        RECT  0.635 1.755 0.895 2.015 ;
        RECT  0.125 0.650 0.385 1.060 ;
    END
END AOI2B1X4MTH

MACRO AOI2B1X8MTH
    CLASS CORE ;
    FOREIGN AOI2B1X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 0.405 6.745 2.085 ;
        RECT  6.155 0.800 6.485 2.085 ;
        RECT  5.725 0.800 6.155 1.070 ;
        RECT  5.440 1.765 6.155 2.085 ;
        RECT  5.465 0.405 5.725 1.070 ;
        RECT  5.455 0.540 5.465 1.070 ;
        RECT  2.130 0.540 5.455 0.810 ;
        END
        AntennaDiffArea 1.884 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.305 1.255 5.935 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.180 0.555 1.505 ;
        RECT  0.100 1.180 0.310 1.735 ;
        END
        AntennaGateArea 0.2054 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.835 0.990 4.435 1.345 ;
        RECT  2.405 0.990 3.835 1.150 ;
        RECT  1.950 0.990 2.405 1.345 ;
        RECT  1.740 0.875 1.950 1.345 ;
        END
        AntennaGateArea 0.8216 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.255 -0.130 7.380 0.130 ;
        RECT  6.995 -0.130 7.255 0.955 ;
        RECT  6.235 -0.130 6.995 0.130 ;
        RECT  5.975 -0.130 6.235 0.620 ;
        RECT  5.155 -0.130 5.975 0.130 ;
        RECT  4.895 -0.130 5.155 0.355 ;
        RECT  3.280 -0.130 4.895 0.130 ;
        RECT  3.020 -0.130 3.280 0.350 ;
        RECT  1.320 -0.130 3.020 0.130 ;
        RECT  0.720 -0.130 1.320 0.650 ;
        RECT  0.000 -0.130 0.720 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.705 2.740 7.380 3.000 ;
        RECT  4.445 2.205 4.705 3.000 ;
        RECT  2.745 2.740 4.445 3.000 ;
        RECT  2.485 2.205 2.745 3.000 ;
        RECT  0.385 2.740 2.485 3.000 ;
        RECT  0.125 1.915 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.995 1.865 7.255 2.465 ;
        RECT  5.215 2.305 6.995 2.465 ;
        RECT  4.955 1.865 5.215 2.465 ;
        RECT  4.195 1.865 4.955 2.025 ;
        RECT  4.665 1.315 4.925 1.685 ;
        RECT  3.425 1.525 4.665 1.685 ;
        RECT  3.935 1.865 4.195 2.465 ;
        RECT  3.255 1.865 3.935 2.025 ;
        RECT  2.805 1.360 3.425 1.685 ;
        RECT  2.995 1.865 3.255 2.465 ;
        RECT  2.235 1.865 2.995 2.025 ;
        RECT  1.545 1.525 2.805 1.685 ;
        RECT  1.975 1.865 2.235 2.490 ;
        RECT  1.295 1.865 1.975 2.025 ;
        RECT  1.285 0.830 1.545 1.685 ;
        RECT  1.135 1.865 1.295 2.515 ;
        RECT  0.385 0.830 1.285 0.990 ;
        RECT  0.895 1.525 1.285 1.685 ;
        RECT  1.035 2.255 1.135 2.515 ;
        RECT  0.735 1.525 0.895 1.945 ;
        RECT  0.635 1.685 0.735 1.945 ;
        RECT  0.125 0.370 0.385 0.990 ;
    END
END AOI2B1X8MTH

MACRO AOI2B1XLMTH
    CLASS CORE ;
    FOREIGN AOI2B1XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.770 2.370 2.025 ;
        RECT  1.540 0.770 2.210 0.930 ;
        RECT  2.125 1.700 2.210 2.025 ;
        END
        AntennaDiffArea 0.25 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.110 2.030 1.460 ;
        RECT  1.730 1.110 1.950 1.585 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.430 1.155 0.730 1.585 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.110 1.550 1.585 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 -0.130 2.460 0.130 ;
        RECT  2.070 -0.130 2.330 0.390 ;
        RECT  1.640 -0.130 2.070 0.130 ;
        RECT  0.700 -0.130 1.640 0.380 ;
        RECT  0.425 -0.130 0.700 0.130 ;
        RECT  0.165 -0.130 0.425 0.390 ;
        RECT  0.000 -0.130 0.165 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 2.740 2.460 3.000 ;
        RECT  1.580 2.305 2.180 3.000 ;
        RECT  1.295 2.740 1.580 3.000 ;
        RECT  0.695 2.305 1.295 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.555 1.770 1.825 1.930 ;
        RECT  0.910 0.815 1.070 1.505 ;
        RECT  0.250 0.815 0.910 0.975 ;
        RECT  0.250 2.355 0.385 2.515 ;
        RECT  0.090 0.815 0.250 2.515 ;
    END
END AOI2B1XLMTH

MACRO AOI2BB1X1MTH
    CLASS CORE ;
    FOREIGN AOI2BB1X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.790 2.370 2.125 ;
        RECT  1.540 0.790 2.210 0.950 ;
        RECT  2.125 1.700 2.210 2.125 ;
        END
        AntennaDiffArea 0.4 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.130 1.605 1.675 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.170 1.130 1.680 ;
        END
        AntennaGateArea 0.065 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.790 0.355 1.475 ;
        END
        AntennaGateArea 0.065 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 -0.130 2.460 0.130 ;
        RECT  1.720 -0.130 2.320 0.390 ;
        RECT  1.175 -0.130 1.720 0.130 ;
        RECT  0.235 -0.130 1.175 0.510 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.310 2.740 2.460 3.000 ;
        RECT  1.710 2.570 2.310 3.000 ;
        RECT  1.285 2.740 1.710 3.000 ;
        RECT  1.025 2.205 1.285 3.000 ;
        RECT  0.750 2.740 1.025 3.000 ;
        RECT  0.150 2.570 0.750 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.945 1.235 2.030 1.495 ;
        RECT  1.785 1.235 1.945 2.025 ;
        RECT  0.695 1.865 1.785 2.025 ;
        RECT  0.695 0.815 0.815 0.975 ;
        RECT  0.535 0.815 0.695 2.025 ;
        RECT  0.125 1.735 0.535 2.025 ;
    END
END AOI2BB1X1MTH

MACRO AOI2BB1X2MTH
    CLASS CORE ;
    FOREIGN AOI2BB1X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.290 1.285 2.360 2.465 ;
        RECT  2.130 0.560 2.290 2.465 ;
        RECT  1.750 0.560 2.130 0.720 ;
        RECT  1.910 2.205 2.130 2.465 ;
        RECT  1.490 0.460 1.750 0.720 ;
        END
        AntennaDiffArea 0.57 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.245 1.605 1.675 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.655 1.245 1.130 1.670 ;
        END
        AntennaGateArea 0.1053 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.980 0.355 1.680 ;
        END
        AntennaGateArea 0.1053 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.290 -0.130 2.460 0.130 ;
        RECT  2.030 -0.130 2.290 0.380 ;
        RECT  1.195 -0.130 2.030 0.130 ;
        RECT  0.205 -0.130 1.195 0.475 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 2.740 2.460 3.000 ;
        RECT  1.015 2.205 1.275 3.000 ;
        RECT  0.785 2.740 1.015 3.000 ;
        RECT  0.185 2.570 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.790 0.905 1.950 2.025 ;
        RECT  0.740 0.905 1.790 1.065 ;
        RECT  0.385 1.865 1.790 2.025 ;
        RECT  0.580 0.765 0.740 1.065 ;
        RECT  0.125 1.865 0.385 2.125 ;
    END
END AOI2BB1X2MTH

MACRO AOI2BB1X4MTH
    CLASS CORE ;
    FOREIGN AOI2BB1X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.880 3.590 2.050 ;
        RECT  3.015 0.880 3.380 1.060 ;
        RECT  2.355 1.870 3.380 2.050 ;
        RECT  2.755 0.385 3.015 1.060 ;
        RECT  1.935 0.540 2.755 0.720 ;
        RECT  2.095 1.870 2.355 2.510 ;
        RECT  1.675 0.460 1.935 0.720 ;
        END
        AntennaDiffArea 1.104 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 1.245 3.155 1.690 ;
        RECT  1.560 1.530 2.895 1.690 ;
        RECT  1.330 1.245 1.560 1.690 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.245 1.150 1.710 ;
        END
        AntennaGateArea 0.1924 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.980 0.355 1.580 ;
        END
        AntennaGateArea 0.1924 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.700 ;
        RECT  2.475 -0.130 3.305 0.130 ;
        RECT  2.215 -0.130 2.475 0.360 ;
        RECT  1.415 -0.130 2.215 0.130 ;
        RECT  1.155 -0.130 1.415 0.715 ;
        RECT  0.385 -0.130 1.155 0.130 ;
        RECT  0.125 -0.130 0.385 0.715 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.365 2.740 3.690 3.000 ;
        RECT  3.105 2.230 3.365 3.000 ;
        RECT  1.315 2.740 3.105 3.000 ;
        RECT  1.055 1.890 1.315 3.000 ;
        RECT  0.000 2.740 1.055 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.040 1.190 2.480 1.350 ;
        RECT  1.880 0.900 2.040 1.350 ;
        RECT  0.895 0.900 1.880 1.060 ;
        RECT  0.695 0.640 0.895 1.060 ;
        RECT  0.635 0.640 0.695 1.995 ;
        RECT  0.535 0.900 0.635 1.995 ;
        RECT  0.385 1.835 0.535 1.995 ;
        RECT  0.125 1.835 0.385 2.435 ;
    END
END AOI2BB1X4MTH

MACRO AOI2BB1X8MTH
    CLASS CORE ;
    FOREIGN AOI2BB1X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.175 0.460 6.460 2.130 ;
        RECT  2.615 0.460 6.175 0.720 ;
        RECT  5.315 1.870 6.175 2.130 ;
        RECT  5.055 1.870 5.315 2.475 ;
        RECT  3.275 1.870 5.055 2.130 ;
        RECT  3.015 1.870 3.275 2.470 ;
        END
        AntennaDiffArea 2.002 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.815 1.205 5.975 1.690 ;
        RECT  4.385 1.530 5.815 1.690 ;
        RECT  3.785 1.245 4.385 1.690 ;
        RECT  2.485 1.530 3.785 1.690 ;
        RECT  2.150 1.245 2.485 1.690 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.830 1.245 1.970 1.580 ;
        RECT  1.670 1.245 1.830 1.885 ;
        RECT  0.605 1.725 1.670 1.885 ;
        RECT  0.445 1.245 0.605 1.885 ;
        END
        AntennaGateArea 0.3848 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.240 1.490 1.540 ;
        END
        AntennaGateArea 0.3848 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.280 ;
        RECT  4.355 -0.130 6.175 0.130 ;
        RECT  4.095 -0.130 4.355 0.270 ;
        RECT  2.355 -0.130 4.095 0.130 ;
        RECT  2.095 -0.130 2.355 0.715 ;
        RECT  0.385 -0.130 2.095 0.130 ;
        RECT  0.125 -0.130 0.385 0.715 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.235 2.740 6.560 3.000 ;
        RECT  5.975 2.310 6.235 3.000 ;
        RECT  4.255 2.740 5.975 3.000 ;
        RECT  3.995 2.315 4.255 3.000 ;
        RECT  2.270 2.740 3.995 3.000 ;
        RECT  2.010 1.925 2.270 3.000 ;
        RECT  0.445 2.740 2.010 3.000 ;
        RECT  0.185 2.405 0.445 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.025 1.095 5.465 1.350 ;
        RECT  4.865 0.900 5.025 1.350 ;
        RECT  3.440 0.900 4.865 1.060 ;
        RECT  2.840 0.900 3.440 1.350 ;
        RECT  1.835 0.900 2.840 1.060 ;
        RECT  1.575 0.640 1.835 1.060 ;
        RECT  0.905 0.900 1.575 1.060 ;
        RECT  1.060 2.065 1.320 2.325 ;
        RECT  0.265 2.065 1.060 2.225 ;
        RECT  0.645 0.640 0.905 1.060 ;
        RECT  0.265 0.900 0.645 1.060 ;
        RECT  0.105 0.900 0.265 2.225 ;
    END
END AOI2BB1X8MTH

MACRO AOI2BB1XLMTH
    CLASS CORE ;
    FOREIGN AOI2BB1XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.310 1.285 2.360 2.030 ;
        RECT  2.150 0.565 2.310 2.030 ;
        RECT  1.555 0.565 2.150 0.725 ;
        RECT  2.110 1.770 2.150 2.030 ;
        END
        AntennaDiffArea 0.368 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.245 1.590 1.700 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.245 1.130 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.980 0.420 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 -0.130 2.460 0.130 ;
        RECT  2.065 -0.130 2.325 0.365 ;
        RECT  1.175 -0.130 2.065 0.130 ;
        RECT  0.235 -0.130 1.175 0.510 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 2.740 2.460 3.000 ;
        RECT  1.575 2.570 2.175 3.000 ;
        RECT  1.285 2.740 1.575 3.000 ;
        RECT  1.025 2.225 1.285 3.000 ;
        RECT  0.775 2.740 1.025 3.000 ;
        RECT  0.175 2.570 0.775 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.950 1.235 1.970 1.495 ;
        RECT  1.930 0.905 1.950 1.495 ;
        RECT  1.770 0.905 1.930 2.040 ;
        RECT  0.765 0.905 1.770 1.065 ;
        RECT  0.385 1.880 1.770 2.040 ;
        RECT  0.605 0.765 0.765 1.065 ;
        RECT  0.125 1.760 0.385 2.040 ;
    END
END AOI2BB1XLMTH

MACRO AOI2BB2X1MTH
    CLASS CORE ;
    FOREIGN AOI2BB2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 1.285 3.180 2.015 ;
        RECT  2.945 0.475 3.130 2.015 ;
        RECT  2.255 0.475 2.945 0.635 ;
        END
        AntennaDiffArea 0.453 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.155 1.785 1.695 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.245 2.425 1.695 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.980 0.355 1.580 ;
        END
        AntennaGateArea 0.065 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.155 1.150 1.700 ;
        END
        AntennaGateArea 0.065 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 -0.130 3.280 0.130 ;
        RECT  2.825 -0.130 3.085 0.295 ;
        RECT  1.620 -0.130 2.825 0.130 ;
        RECT  1.360 -0.130 1.620 0.590 ;
        RECT  1.065 -0.130 1.360 0.130 ;
        RECT  0.125 -0.130 1.065 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 2.740 3.280 3.000 ;
        RECT  2.465 2.570 3.065 3.000 ;
        RECT  2.095 2.740 2.465 3.000 ;
        RECT  1.155 2.555 2.095 3.000 ;
        RECT  0.725 2.740 1.155 3.000 ;
        RECT  0.125 2.380 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.605 0.815 2.765 1.495 ;
        RECT  1.400 1.880 2.645 2.040 ;
        RECT  0.695 0.815 2.605 0.975 ;
        RECT  0.695 1.880 1.145 2.040 ;
        RECT  0.535 0.815 0.695 2.040 ;
    END
END AOI2BB2X1MTH

MACRO AOI2BB2X2MTH
    CLASS CORE ;
    FOREIGN AOI2BB2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 1.290 3.180 2.355 ;
        RECT  2.905 0.475 3.125 2.355 ;
        RECT  2.390 0.475 2.905 0.635 ;
        RECT  2.855 1.755 2.905 2.355 ;
        RECT  2.130 0.375 2.390 0.635 ;
        END
        AntennaDiffArea 0.636 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.155 1.770 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.155 2.360 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.980 0.355 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.155 1.150 1.625 ;
        END
        AntennaGateArea 0.1053 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.985 -0.130 3.280 0.130 ;
        RECT  2.725 -0.130 2.985 0.295 ;
        RECT  1.420 -0.130 2.725 0.130 ;
        RECT  1.160 -0.130 1.420 0.590 ;
        RECT  0.725 -0.130 1.160 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 2.740 3.280 3.000 ;
        RECT  1.795 2.110 2.055 3.000 ;
        RECT  0.730 2.740 1.795 3.000 ;
        RECT  0.130 2.450 0.730 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.565 0.815 2.725 1.495 ;
        RECT  2.345 1.770 2.605 2.390 ;
        RECT  0.695 0.815 2.565 0.975 ;
        RECT  1.525 1.770 2.345 1.930 ;
        RECT  1.365 1.770 1.525 2.515 ;
        RECT  1.245 2.255 1.365 2.515 ;
        RECT  0.695 1.805 1.105 1.965 ;
        RECT  0.535 0.815 0.695 1.965 ;
    END
END AOI2BB2X2MTH

MACRO AOI2BB2X4MTH
    CLASS CORE ;
    FOREIGN AOI2BB2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.470 0.550 3.730 0.810 ;
        RECT  2.215 0.630 3.470 0.810 ;
        RECT  2.215 1.245 2.360 1.585 ;
        RECT  2.015 0.375 2.215 2.115 ;
        RECT  1.905 0.375 2.015 0.975 ;
        RECT  1.905 1.855 2.015 2.115 ;
        END
        AntennaDiffArea 0.876 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.135 0.990 4.395 1.495 ;
        RECT  3.035 0.990 4.135 1.150 ;
        RECT  2.560 0.990 3.035 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.285 1.330 3.900 1.585 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.255 0.645 1.580 ;
        END
        AntennaGateArea 0.1924 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.245 1.380 1.580 ;
        END
        AntennaGateArea 0.1924 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.605 -0.130 4.920 0.130 ;
        RECT  4.345 -0.130 4.605 0.730 ;
        RECT  2.790 -0.130 4.345 0.130 ;
        RECT  2.530 -0.130 2.790 0.445 ;
        RECT  1.545 -0.130 2.530 0.130 ;
        RECT  1.285 -0.130 1.545 0.640 ;
        RECT  0.385 -0.130 1.285 0.130 ;
        RECT  0.125 -0.130 0.385 0.755 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.255 2.740 4.920 3.000 ;
        RECT  3.995 2.135 4.255 3.000 ;
        RECT  3.215 2.740 3.995 3.000 ;
        RECT  2.955 2.165 3.215 3.000 ;
        RECT  0.385 2.740 2.955 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.510 1.765 4.770 2.365 ;
        RECT  3.735 1.765 4.510 1.925 ;
        RECT  3.475 1.765 3.735 2.435 ;
        RECT  2.695 1.765 3.475 1.925 ;
        RECT  2.435 1.765 2.695 2.525 ;
        RECT  1.655 2.365 2.435 2.525 ;
        RECT  1.720 1.245 1.835 1.505 ;
        RECT  1.560 0.900 1.720 1.920 ;
        RECT  1.395 2.255 1.655 2.525 ;
        RECT  0.905 0.900 1.560 1.060 ;
        RECT  0.955 1.760 1.560 1.920 ;
        RECT  0.645 0.645 0.905 1.060 ;
    END
END AOI2BB2X4MTH

MACRO AOI2BB2X8MTH
    CLASS CORE ;
    FOREIGN AOI2BB2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.105 0.480 7.465 0.770 ;
        RECT  4.075 0.480 4.105 1.055 ;
        RECT  4.040 0.375 4.075 1.055 ;
        RECT  3.815 0.375 4.040 2.195 ;
        RECT  3.775 0.775 3.815 2.195 ;
        RECT  3.380 0.775 3.775 2.075 ;
        RECT  2.995 0.775 3.380 1.055 ;
        RECT  2.735 1.725 3.380 2.075 ;
        RECT  2.735 0.375 2.995 1.055 ;
        END
        AntennaDiffArea 1.914 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.955 1.205 8.195 1.465 ;
        RECT  7.795 0.990 7.955 1.465 ;
        RECT  6.620 0.990 7.795 1.150 ;
        RECT  6.020 0.990 6.620 1.345 ;
        RECT  4.835 0.990 6.020 1.150 ;
        RECT  4.410 0.990 4.835 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.965 1.330 7.565 1.685 ;
        RECT  5.695 1.525 6.965 1.685 ;
        RECT  5.055 1.330 5.695 1.685 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.775 1.290 1.375 1.580 ;
        END
        AntennaGateArea 0.3848 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.570 0.950 2.050 1.580 ;
        RECT  0.555 0.950 1.570 1.110 ;
        RECT  0.295 0.950 0.555 1.505 ;
        END
        AntennaGateArea 0.3848 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.405 -0.130 8.610 0.130 ;
        RECT  8.145 -0.130 8.405 0.980 ;
        RECT  6.480 -0.130 8.145 0.130 ;
        RECT  6.220 -0.130 6.480 0.300 ;
        RECT  4.620 -0.130 6.220 0.130 ;
        RECT  4.360 -0.130 4.620 0.300 ;
        RECT  3.535 -0.130 4.360 0.130 ;
        RECT  3.275 -0.130 3.535 0.590 ;
        RECT  2.455 -0.130 3.275 0.130 ;
        RECT  2.195 -0.130 2.455 0.430 ;
        RECT  0.385 -0.130 2.195 0.130 ;
        RECT  0.125 -0.130 0.385 0.770 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.965 2.740 8.610 3.000 ;
        RECT  7.705 2.205 7.965 3.000 ;
        RECT  5.065 2.740 7.705 3.000 ;
        RECT  4.805 2.205 5.065 3.000 ;
        RECT  1.215 2.740 4.805 3.000 ;
        RECT  0.955 2.150 1.215 3.000 ;
        RECT  0.000 2.740 0.955 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.225 1.865 8.485 2.465 ;
        RECT  7.455 1.865 8.225 2.025 ;
        RECT  7.195 1.865 7.455 2.480 ;
        RECT  6.515 1.865 7.195 2.025 ;
        RECT  6.255 1.865 6.515 2.475 ;
        RECT  5.575 1.865 6.255 2.025 ;
        RECT  5.315 1.865 5.575 2.475 ;
        RECT  4.545 1.865 5.315 2.025 ;
        RECT  4.285 1.865 4.545 2.560 ;
        RECT  3.525 2.400 4.285 2.560 ;
        RECT  3.265 2.255 3.525 2.560 ;
        RECT  2.485 2.400 3.265 2.560 ;
        RECT  2.550 1.245 3.155 1.505 ;
        RECT  2.390 0.610 2.550 1.920 ;
        RECT  2.225 2.255 2.485 2.560 ;
        RECT  1.915 0.610 2.390 0.770 ;
        RECT  0.385 1.760 2.390 1.920 ;
        RECT  1.655 0.510 1.915 0.770 ;
        RECT  0.895 0.610 1.655 0.770 ;
        RECT  0.635 0.510 0.895 0.770 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END AOI2BB2X8MTH

MACRO AOI2BB2XLMTH
    CLASS CORE ;
    FOREIGN AOI2BB2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.645 1.695 2.770 2.035 ;
        RECT  2.485 0.815 2.645 2.035 ;
        RECT  1.985 0.815 2.485 0.975 ;
        END
        AntennaDiffArea 0.238 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.060 1.560 1.900 ;
        END
        AntennaGateArea 0.0663 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.170 2.285 1.620 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.865 0.350 1.705 ;
        END
        AntennaGateArea 0.0624 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 1.045 1.150 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 2.870 0.130 ;
        RECT  2.485 -0.130 2.745 0.250 ;
        RECT  1.215 -0.130 2.485 0.130 ;
        RECT  0.275 -0.130 1.215 0.385 ;
        RECT  0.000 -0.130 0.275 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.735 2.740 2.870 3.000 ;
        RECT  2.475 2.570 2.735 3.000 ;
        RECT  2.165 2.740 2.475 3.000 ;
        RECT  1.565 2.445 2.165 3.000 ;
        RECT  0.725 2.740 1.565 3.000 ;
        RECT  0.125 2.265 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.805 0.445 2.365 0.605 ;
        RECT  1.975 1.815 2.235 2.260 ;
        RECT  1.275 2.100 1.975 2.260 ;
        RECT  1.645 0.445 1.805 0.865 ;
        RECT  0.690 0.705 1.645 0.865 ;
        RECT  1.015 2.100 1.275 2.480 ;
        RECT  0.690 1.760 1.145 1.920 ;
        RECT  0.530 0.705 0.690 1.920 ;
    END
END AOI2BB2XLMTH

MACRO AOI31X1MTH
    CLASS CORE ;
    FOREIGN AOI31X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.770 2.370 2.085 ;
        RECT  1.510 0.770 2.210 0.930 ;
        RECT  2.150 1.700 2.210 2.085 ;
        RECT  2.125 1.825 2.150 2.085 ;
        END
        AntennaDiffArea 0.363 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.115 2.030 1.465 ;
        RECT  1.740 1.115 1.950 1.665 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.325 1.350 0.640 1.665 ;
        RECT  0.100 1.290 0.325 1.665 ;
        END
        AntennaGateArea 0.1274 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 0.880 1.100 1.485 ;
        RECT  0.510 0.880 0.840 1.170 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 1.110 1.550 1.665 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 -0.130 2.460 0.130 ;
        RECT  2.070 -0.130 2.330 0.590 ;
        RECT  1.720 -0.130 2.070 0.130 ;
        RECT  0.780 -0.130 1.720 0.385 ;
        RECT  0.415 -0.130 0.780 0.130 ;
        RECT  0.155 -0.130 0.415 0.685 ;
        RECT  0.000 -0.130 0.155 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 2.740 2.460 3.000 ;
        RECT  1.445 2.555 2.045 3.000 ;
        RECT  1.170 2.740 1.445 3.000 ;
        RECT  0.230 2.555 1.170 3.000 ;
        RECT  0.000 2.740 0.230 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.565 1.845 1.825 2.065 ;
    END
END AOI31X1MTH

MACRO AOI31X2MTH
    CLASS CORE ;
    FOREIGN AOI31X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.770 2.370 2.430 ;
        RECT  1.740 0.770 2.210 0.930 ;
        RECT  2.075 1.830 2.210 2.430 ;
        RECT  1.480 0.405 1.740 0.930 ;
        END
        AntennaDiffArea 0.566 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 1.115 2.030 1.465 ;
        RECT  1.740 1.115 1.970 1.670 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.325 1.365 0.640 1.685 ;
        RECT  0.100 1.290 0.325 1.685 ;
        END
        AntennaGateArea 0.2054 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.820 0.880 1.070 1.485 ;
        RECT  0.510 0.880 0.820 1.170 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.110 1.550 1.695 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.310 -0.130 2.460 0.130 ;
        RECT  2.050 -0.130 2.310 0.590 ;
        RECT  0.385 -0.130 2.050 0.130 ;
        RECT  0.125 -0.130 0.385 0.660 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 2.740 2.460 3.000 ;
        RECT  1.055 2.255 1.315 3.000 ;
        RECT  0.000 2.740 1.055 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.565 1.875 1.825 2.475 ;
        RECT  0.795 1.875 1.565 2.035 ;
        RECT  0.535 1.875 0.795 2.475 ;
    END
END AOI31X2MTH

MACRO AOI31X4MTH
    CLASS CORE ;
    FOREIGN AOI31X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.320 0.380 4.570 1.170 ;
        RECT  4.310 0.380 4.320 2.160 ;
        RECT  4.090 0.880 4.310 2.160 ;
        RECT  3.455 0.880 4.090 1.060 ;
        RECT  3.940 1.900 4.090 2.160 ;
        RECT  3.195 0.385 3.455 1.060 ;
        RECT  0.660 0.545 3.195 0.725 ;
        RECT  0.400 0.405 0.660 1.005 ;
        END
        AntennaDiffArea 1.132 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 1.255 3.885 1.665 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.580 1.245 2.210 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.670 1.215 2.770 1.475 ;
        RECT  2.510 0.905 2.670 1.475 ;
        RECT  1.310 0.905 2.510 1.065 ;
        RECT  0.880 0.905 1.310 1.485 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 1.240 3.200 1.880 ;
        RECT  0.675 1.720 3.040 1.880 ;
        RECT  0.515 1.225 0.675 1.880 ;
        RECT  0.100 1.225 0.515 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.030 -0.130 4.920 0.130 ;
        RECT  3.770 -0.130 4.030 0.700 ;
        RECT  2.020 -0.130 3.770 0.130 ;
        RECT  1.760 -0.130 2.020 0.365 ;
        RECT  0.000 -0.130 1.760 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.140 2.740 4.920 3.000 ;
        RECT  2.880 2.410 3.140 3.000 ;
        RECT  2.040 2.740 2.880 3.000 ;
        RECT  1.780 2.405 2.040 3.000 ;
        RECT  0.935 2.740 1.780 3.000 ;
        RECT  0.675 2.410 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.500 1.810 4.710 2.520 ;
        RECT  3.690 2.360 4.500 2.520 ;
        RECT  3.430 1.900 3.690 2.520 ;
        RECT  2.590 2.060 3.430 2.220 ;
        RECT  2.330 2.060 2.590 2.320 ;
        RECT  1.490 2.060 2.330 2.220 ;
        RECT  1.230 2.060 1.490 2.320 ;
        RECT  0.385 2.060 1.230 2.220 ;
        RECT  0.125 2.060 0.385 2.320 ;
    END
END AOI31X4MTH

MACRO AOI31XLMTH
    CLASS CORE ;
    FOREIGN AOI31XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.770 2.370 2.085 ;
        RECT  1.540 0.770 2.210 0.930 ;
        RECT  2.150 1.700 2.210 2.085 ;
        RECT  2.125 1.825 2.150 2.085 ;
        END
        AntennaDiffArea 0.25 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 1.115 2.030 1.465 ;
        RECT  1.740 1.115 1.970 1.685 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.325 1.365 0.640 1.685 ;
        RECT  0.100 1.290 0.325 1.685 ;
        END
        AntennaGateArea 0.0702 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.820 0.880 1.120 1.505 ;
        RECT  0.510 0.880 0.820 1.170 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 1.110 1.550 1.695 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  2.075 -0.130 2.335 0.470 ;
        RECT  1.720 -0.130 2.075 0.130 ;
        RECT  0.780 -0.130 1.720 0.385 ;
        RECT  0.430 -0.130 0.780 0.130 ;
        RECT  0.170 -0.130 0.430 0.685 ;
        RECT  0.000 -0.130 0.170 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 2.740 2.460 3.000 ;
        RECT  1.630 2.570 2.230 3.000 ;
        RECT  1.170 2.740 1.630 3.000 ;
        RECT  0.230 2.375 1.170 3.000 ;
        RECT  0.000 2.740 0.230 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.565 1.875 1.825 2.035 ;
    END
END AOI31XLMTH

MACRO AOI32X1MTH
    CLASS CORE ;
    FOREIGN AOI32X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.290 0.770 2.400 1.130 ;
        RECT  2.130 0.770 2.290 2.035 ;
        RECT  2.110 0.770 2.130 1.130 ;
        RECT  1.975 1.875 2.130 2.035 ;
        RECT  1.560 0.770 2.110 0.930 ;
        END
        AntennaDiffArea 0.422 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.580 1.005 2.770 1.635 ;
        RECT  2.560 1.290 2.580 1.635 ;
        RECT  2.470 1.310 2.560 1.635 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.650 1.225 1.950 1.695 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.315 0.355 1.985 ;
        RECT  0.100 1.290 0.310 1.985 ;
        END
        AntennaGateArea 0.1274 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.365 1.040 1.525 ;
        RECT  0.560 0.880 0.720 1.525 ;
        RECT  0.510 0.880 0.560 1.170 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.380 1.225 1.470 1.485 ;
        RECT  1.220 0.880 1.380 1.485 ;
        RECT  0.920 0.880 1.220 1.170 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 2.870 0.130 ;
        RECT  2.485 -0.130 2.745 0.590 ;
        RECT  2.245 -0.130 2.485 0.130 ;
        RECT  1.305 -0.130 2.245 0.385 ;
        RECT  1.065 -0.130 1.305 0.130 ;
        RECT  0.125 -0.130 1.065 0.385 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.535 2.740 2.870 3.000 ;
        RECT  1.595 2.555 2.535 3.000 ;
        RECT  1.170 2.740 1.595 3.000 ;
        RECT  0.230 2.555 1.170 3.000 ;
        RECT  0.000 2.740 0.230 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.535 1.825 2.695 2.375 ;
        RECT  1.725 2.215 2.535 2.375 ;
        RECT  1.465 1.890 1.725 2.375 ;
        RECT  0.535 1.890 1.465 2.150 ;
    END
END AOI32X1MTH

MACRO AOI32X2MTH
    CLASS CORE ;
    FOREIGN AOI32X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.785 3.180 2.010 ;
        RECT  1.985 0.785 2.970 0.945 ;
        RECT  2.585 1.850 2.970 2.010 ;
        RECT  2.325 1.850 2.585 2.110 ;
        RECT  1.725 0.440 1.985 0.945 ;
        END
        AntennaDiffArea 0.77 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.540 1.125 2.790 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 1.125 2.360 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.345 1.065 0.720 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.955 1.150 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.125 1.735 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 -0.130 3.280 0.130 ;
        RECT  2.675 -0.130 2.935 0.590 ;
        RECT  0.510 -0.130 2.675 0.130 ;
        RECT  0.250 -0.130 0.510 0.745 ;
        RECT  0.000 -0.130 0.250 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.525 2.740 3.280 3.000 ;
        RECT  1.265 2.100 1.525 3.000 ;
        RECT  0.425 2.740 1.265 3.000 ;
        RECT  0.165 1.805 0.425 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.845 2.190 3.105 2.460 ;
        RECT  2.075 2.300 2.845 2.460 ;
        RECT  1.815 1.760 2.075 2.460 ;
        RECT  0.975 1.760 1.815 1.920 ;
        RECT  0.715 1.760 0.975 2.365 ;
    END
END AOI32X2MTH

MACRO AOI32X4MTH
    CLASS CORE ;
    FOREIGN AOI32X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.430 0.385 5.640 2.080 ;
        RECT  5.210 0.385 5.430 0.985 ;
        RECT  3.795 1.900 5.430 2.080 ;
        RECT  3.755 0.540 5.210 0.740 ;
        RECT  3.155 0.355 3.755 0.955 ;
        RECT  0.395 0.550 3.155 0.810 ;
        RECT  0.135 0.370 0.395 0.970 ;
        END
        AntennaDiffArea 1.662 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.180 0.920 4.860 1.380 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.090 1.310 5.250 1.720 ;
        RECT  4.000 1.560 5.090 1.720 ;
        RECT  3.685 1.210 4.000 1.720 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.515 1.330 2.180 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 0.990 2.810 1.540 ;
        RECT  1.095 0.990 2.360 1.150 ;
        RECT  0.935 0.990 1.095 1.520 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.150 1.225 3.270 1.485 ;
        RECT  2.990 1.225 3.150 1.880 ;
        RECT  0.660 1.720 2.990 1.880 ;
        RECT  0.500 1.225 0.660 1.880 ;
        RECT  0.100 1.225 0.500 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.615 -0.130 5.740 0.130 ;
        RECT  4.355 -0.130 4.615 0.360 ;
        RECT  1.955 -0.130 4.355 0.130 ;
        RECT  1.695 -0.130 1.955 0.365 ;
        RECT  0.000 -0.130 1.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.005 2.740 5.740 3.000 ;
        RECT  2.745 2.405 3.005 3.000 ;
        RECT  0.935 2.740 2.745 3.000 ;
        RECT  0.675 2.435 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.505 2.260 5.615 2.420 ;
        RECT  3.345 1.775 3.505 2.420 ;
        RECT  2.455 2.060 3.345 2.220 ;
        RECT  2.195 2.060 2.455 2.320 ;
        RECT  1.485 2.060 2.195 2.220 ;
        RECT  1.225 2.060 1.485 2.320 ;
        RECT  0.385 2.060 1.225 2.220 ;
        RECT  0.125 2.060 0.385 2.320 ;
    END
END AOI32X4MTH

MACRO AOI32XLMTH
    CLASS CORE ;
    FOREIGN AOI32XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.290 0.820 2.400 1.130 ;
        RECT  2.130 0.720 2.290 1.970 ;
        RECT  2.110 0.720 2.130 1.130 ;
        RECT  2.125 1.710 2.130 1.970 ;
        RECT  1.600 0.720 2.110 0.980 ;
        END
        AntennaDiffArea 0.288 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.290 2.770 1.895 ;
        RECT  2.470 1.315 2.560 1.895 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.940 1.290 1.950 1.580 ;
        RECT  1.890 1.290 1.940 1.695 ;
        RECT  1.650 1.160 1.890 1.695 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.315 0.355 1.685 ;
        RECT  0.100 1.025 0.310 1.685 ;
        END
        AntennaGateArea 0.0702 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.365 1.040 1.525 ;
        RECT  0.560 0.880 0.720 1.525 ;
        RECT  0.510 0.880 0.560 1.170 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.415 1.225 1.470 1.485 ;
        RECT  1.255 0.880 1.415 1.485 ;
        RECT  0.920 0.880 1.255 1.170 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 2.870 0.130 ;
        RECT  2.485 -0.130 2.745 0.590 ;
        RECT  2.245 -0.130 2.485 0.130 ;
        RECT  1.305 -0.130 2.245 0.385 ;
        RECT  1.065 -0.130 1.305 0.130 ;
        RECT  0.125 -0.130 1.065 0.385 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.170 2.740 2.870 3.000 ;
        RECT  0.230 2.375 1.170 3.000 ;
        RECT  0.000 2.740 0.230 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.750 2.295 2.615 2.555 ;
        RECT  1.590 1.875 1.750 2.555 ;
        RECT  0.860 1.875 1.590 2.035 ;
        RECT  0.600 1.795 0.860 2.035 ;
    END
END AOI32XLMTH

MACRO AOI33X1MTH
    CLASS CORE ;
    FOREIGN AOI33X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.715 3.590 2.115 ;
        RECT  1.520 0.715 3.380 0.915 ;
        RECT  3.305 1.770 3.380 2.115 ;
        RECT  2.225 1.770 3.305 1.930 ;
        END
        AntennaDiffArea 0.707 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.600 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.780 0.855 1.130 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.100 1.560 1.665 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.095 3.200 1.590 ;
        END
        AntennaGateArea 0.1274 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 1.095 2.770 1.590 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.110 2.240 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 -0.130 3.690 0.130 ;
        RECT  3.200 -0.130 3.460 0.530 ;
        RECT  2.985 -0.130 3.200 0.130 ;
        RECT  2.045 -0.130 2.985 0.390 ;
        RECT  1.660 -0.130 2.045 0.130 ;
        RECT  0.720 -0.130 1.660 0.390 ;
        RECT  0.440 -0.130 0.720 0.130 ;
        RECT  0.180 -0.130 0.440 1.025 ;
        RECT  0.000 -0.130 0.180 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.555 2.740 3.690 3.000 ;
        RECT  2.955 2.570 3.555 3.000 ;
        RECT  2.660 2.740 2.955 3.000 ;
        RECT  1.720 2.570 2.660 3.000 ;
        RECT  1.420 2.740 1.720 3.000 ;
        RECT  0.820 2.570 1.420 3.000 ;
        RECT  0.385 2.740 0.820 3.000 ;
        RECT  0.125 1.865 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.975 2.110 3.025 2.270 ;
        RECT  1.715 1.850 1.975 2.270 ;
        RECT  0.645 1.850 1.715 2.110 ;
    END
END AOI33X1MTH

MACRO AOI33X2MTH
    CLASS CORE ;
    FOREIGN AOI33X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.785 3.590 2.445 ;
        RECT  2.120 0.785 3.380 0.965 ;
        RECT  3.290 1.825 3.380 2.445 ;
        RECT  2.515 1.825 3.290 2.085 ;
        RECT  2.255 1.825 2.515 2.185 ;
        RECT  1.520 0.365 2.120 0.965 ;
        END
        AntennaDiffArea 1.142 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.580 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.770 0.985 1.130 1.660 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.145 1.560 1.660 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.145 3.200 1.640 ;
        END
        AntennaGateArea 0.2054 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.425 1.145 2.770 1.640 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.145 2.240 1.640 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 -0.130 3.690 0.130 ;
        RECT  3.200 -0.130 3.460 0.605 ;
        RECT  0.395 -0.130 3.200 0.130 ;
        RECT  0.135 -0.130 0.395 1.025 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.480 2.740 3.690 3.000 ;
        RECT  1.220 2.205 1.480 3.000 ;
        RECT  0.400 2.740 1.220 3.000 ;
        RECT  0.140 1.835 0.400 3.000 ;
        RECT  0.000 2.740 0.140 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.775 2.265 3.035 2.525 ;
        RECT  2.005 2.365 2.775 2.525 ;
        RECT  1.745 1.840 2.005 2.525 ;
        RECT  0.950 1.840 1.745 2.000 ;
        RECT  0.690 1.840 0.950 2.440 ;
    END
END AOI33X2MTH

MACRO AOI33X4MTH
    CLASS CORE ;
    FOREIGN AOI33X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.685 0.385 6.870 2.150 ;
        RECT  6.660 0.385 6.685 1.170 ;
        RECT  3.805 1.990 6.685 2.150 ;
        RECT  6.465 0.385 6.660 0.985 ;
        RECT  3.520 0.550 6.465 0.730 ;
        RECT  3.260 0.355 3.520 0.955 ;
        RECT  0.395 0.550 3.260 0.730 ;
        RECT  0.135 0.370 0.395 0.970 ;
        END
        AntennaDiffArea 1.842 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.430 1.330 2.230 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 0.990 2.810 1.540 ;
        RECT  1.145 0.990 2.440 1.150 ;
        RECT  0.885 0.990 1.145 1.500 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.035 1.225 3.195 1.880 ;
        RECT  0.565 1.720 3.035 1.880 ;
        RECT  0.100 1.225 0.565 1.880 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.715 0.910 5.575 1.130 ;
        END
        AntennaGateArea 0.4108 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.815 1.210 6.075 1.470 ;
        RECT  4.455 1.310 5.815 1.470 ;
        RECT  3.985 0.920 4.455 1.470 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.345 1.305 6.505 1.810 ;
        RECT  3.675 1.650 6.345 1.810 ;
        RECT  3.380 1.225 3.675 1.810 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.320 -0.130 6.970 0.130 ;
        RECT  4.720 -0.130 5.320 0.365 ;
        RECT  1.965 -0.130 4.720 0.130 ;
        RECT  1.705 -0.130 1.965 0.365 ;
        RECT  0.000 -0.130 1.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.005 2.740 6.970 3.000 ;
        RECT  2.745 2.405 3.005 3.000 ;
        RECT  0.935 2.740 2.745 3.000 ;
        RECT  0.675 2.435 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.555 2.335 6.785 2.495 ;
        RECT  3.295 2.060 3.555 2.495 ;
        RECT  2.455 2.060 3.295 2.220 ;
        RECT  2.195 2.060 2.455 2.320 ;
        RECT  1.485 2.060 2.195 2.220 ;
        RECT  1.225 2.060 1.485 2.320 ;
        RECT  0.385 2.060 1.225 2.220 ;
        RECT  0.125 2.060 0.385 2.320 ;
    END
END AOI33X4MTH

MACRO AOI33XLMTH
    CLASS CORE ;
    FOREIGN AOI33XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.705 3.590 1.975 ;
        RECT  1.670 0.705 3.380 0.965 ;
        RECT  2.165 1.815 3.380 1.975 ;
        END
        AntennaDiffArea 0.486 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.600 1.675 ;
        END
        AntennaGateArea 0.0702 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.780 1.145 1.130 1.695 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.160 1.560 1.695 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.145 3.200 1.635 ;
        END
        AntennaGateArea 0.0702 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 1.145 2.770 1.635 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.145 2.240 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 -0.130 3.690 0.130 ;
        RECT  3.200 -0.130 3.460 0.525 ;
        RECT  2.985 -0.130 3.200 0.130 ;
        RECT  2.045 -0.130 2.985 0.390 ;
        RECT  1.660 -0.130 2.045 0.130 ;
        RECT  0.720 -0.130 1.660 0.390 ;
        RECT  0.440 -0.130 0.720 0.130 ;
        RECT  0.180 -0.130 0.440 1.025 ;
        RECT  0.000 -0.130 0.180 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.530 2.740 3.690 3.000 ;
        RECT  3.270 2.570 3.530 3.000 ;
        RECT  2.230 2.740 3.270 3.000 ;
        RECT  1.630 2.570 2.230 3.000 ;
        RECT  1.205 2.740 1.630 3.000 ;
        RECT  0.265 2.375 1.205 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.915 2.155 2.995 2.315 ;
        RECT  1.755 1.875 1.915 2.315 ;
        RECT  0.585 1.875 1.755 2.035 ;
    END
END AOI33XLMTH

MACRO BUFX10MTH
    CLASS CORE ;
    FOREIGN BUFX10MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.715 0.410 3.975 1.110 ;
        RECT  3.715 1.735 3.975 2.235 ;
        RECT  2.975 0.820 3.715 1.110 ;
        RECT  2.975 1.735 3.715 2.025 ;
        RECT  2.935 0.820 2.975 2.025 ;
        RECT  2.675 0.410 2.935 2.235 ;
        RECT  2.355 0.820 2.675 2.025 ;
        RECT  1.915 0.820 2.355 1.110 ;
        RECT  1.915 1.735 2.355 2.025 ;
        RECT  1.655 0.420 1.915 1.110 ;
        RECT  1.655 1.735 1.915 2.235 ;
        END
        AntennaDiffArea 1.737 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.590 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 -0.130 4.100 0.130 ;
        RECT  3.195 -0.130 3.455 0.640 ;
        RECT  2.425 -0.130 3.195 0.130 ;
        RECT  2.165 -0.130 2.425 0.640 ;
        RECT  1.405 -0.130 2.165 0.130 ;
        RECT  1.145 -0.130 1.405 0.975 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.975 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 2.740 4.100 3.000 ;
        RECT  3.195 2.255 3.455 3.000 ;
        RECT  2.425 2.740 3.195 3.000 ;
        RECT  2.165 2.255 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 1.915 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.830 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.935 1.300 2.085 1.510 ;
        RECT  0.775 0.420 0.935 2.425 ;
        RECT  0.635 0.420 0.775 1.020 ;
        RECT  0.635 1.825 0.775 2.425 ;
    END
END BUFX10MTH

MACRO BUFX12MTH
    CLASS CORE ;
    FOREIGN BUFX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.035 0.595 4.295 1.145 ;
        RECT  4.035 1.655 4.295 2.285 ;
        RECT  3.385 0.745 4.035 1.145 ;
        RECT  3.385 1.655 4.035 2.055 ;
        RECT  3.275 0.745 3.385 2.055 ;
        RECT  3.015 0.420 3.275 2.335 ;
        RECT  2.765 0.555 3.015 2.235 ;
        RECT  2.345 0.555 2.765 1.095 ;
        RECT  2.345 1.695 2.765 2.235 ;
        RECT  2.085 0.420 2.345 1.095 ;
        RECT  2.085 1.695 2.345 2.335 ;
        END
        AntennaDiffArea 1.767 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.290 0.895 1.580 ;
        END
        AntennaGateArea 0.5278 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.795 -0.130 4.920 0.130 ;
        RECT  4.535 -0.130 4.795 0.300 ;
        RECT  3.785 -0.130 4.535 0.130 ;
        RECT  3.525 -0.130 3.785 0.565 ;
        RECT  1.835 -0.130 3.525 0.130 ;
        RECT  1.575 -0.130 1.835 0.975 ;
        RECT  0.785 -0.130 1.575 0.130 ;
        RECT  0.185 -0.130 0.785 0.365 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.795 2.740 4.920 3.000 ;
        RECT  4.535 2.570 4.795 3.000 ;
        RECT  3.785 2.740 4.535 3.000 ;
        RECT  3.525 2.235 3.785 3.000 ;
        RECT  1.835 2.740 3.525 3.000 ;
        RECT  1.575 1.775 1.835 3.000 ;
        RECT  0.785 2.740 1.575 3.000 ;
        RECT  0.185 2.425 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.325 1.315 2.525 1.475 ;
        RECT  1.165 0.420 1.325 2.390 ;
        RECT  1.065 0.420 1.165 1.020 ;
        RECT  1.065 1.790 1.165 2.390 ;
        RECT  0.385 0.860 1.065 1.020 ;
        RECT  0.385 1.790 1.065 1.950 ;
        RECT  0.125 0.760 0.385 1.020 ;
        RECT  0.125 1.790 0.385 2.055 ;
    END
END BUFX12MTH

MACRO BUFX14MTH
    CLASS CORE ;
    FOREIGN BUFX14MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.355 0.425 5.615 2.335 ;
        RECT  4.535 1.085 5.355 1.785 ;
        RECT  4.275 0.425 4.535 2.335 ;
        RECT  3.515 1.085 4.275 1.785 ;
        RECT  3.255 0.420 3.515 2.335 ;
        RECT  2.975 0.745 3.255 2.055 ;
        RECT  2.495 0.745 2.975 1.135 ;
        RECT  2.495 1.655 2.975 2.055 ;
        RECT  2.235 0.420 2.495 1.135 ;
        RECT  2.235 1.655 2.495 2.335 ;
        END
        AntennaDiffArea 2.337 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.290 1.045 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 -0.130 5.740 0.130 ;
        RECT  4.815 -0.130 5.075 0.905 ;
        RECT  4.025 -0.130 4.815 0.130 ;
        RECT  3.765 -0.130 4.025 0.905 ;
        RECT  3.005 -0.130 3.765 0.130 ;
        RECT  2.745 -0.130 3.005 0.565 ;
        RECT  1.985 -0.130 2.745 0.130 ;
        RECT  1.725 -0.130 1.985 0.960 ;
        RECT  0.935 -0.130 1.725 0.130 ;
        RECT  0.675 -0.130 0.935 0.640 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 2.740 5.740 3.000 ;
        RECT  4.815 1.965 5.075 3.000 ;
        RECT  4.025 2.740 4.815 3.000 ;
        RECT  3.765 1.965 4.025 3.000 ;
        RECT  3.005 2.740 3.765 3.000 ;
        RECT  2.745 2.235 3.005 3.000 ;
        RECT  1.985 2.740 2.745 3.000 ;
        RECT  1.725 1.775 1.985 3.000 ;
        RECT  0.935 2.740 1.725 3.000 ;
        RECT  0.675 2.130 0.935 3.000 ;
        RECT  0.000 2.740 0.675 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.475 1.315 2.670 1.475 ;
        RECT  1.315 0.420 1.475 2.390 ;
        RECT  1.215 0.420 1.315 1.020 ;
        RECT  1.215 1.790 1.315 2.390 ;
        RECT  0.395 0.860 1.215 1.020 ;
        RECT  0.395 1.790 1.215 1.950 ;
        RECT  0.135 0.420 0.395 1.020 ;
        RECT  0.135 1.790 0.395 2.390 ;
    END
END BUFX14MTH

MACRO BUFX16MTH
    CLASS CORE ;
    FOREIGN BUFX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.255 0.395 5.515 2.335 ;
        RECT  4.495 1.085 5.255 1.785 ;
        RECT  4.235 0.395 4.495 2.335 ;
        RECT  3.475 1.085 4.235 1.785 ;
        RECT  3.215 0.395 3.475 2.335 ;
        RECT  3.025 0.745 3.215 2.125 ;
        RECT  2.455 0.745 3.025 1.145 ;
        RECT  2.455 1.735 3.025 2.125 ;
        RECT  2.195 0.390 2.455 1.145 ;
        RECT  2.195 1.735 2.455 2.335 ;
        END
        AntennaDiffArea 2.344 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.290 1.065 1.580 ;
        END
        AntennaGateArea 0.6006 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 -0.130 6.150 0.130 ;
        RECT  5.765 -0.130 6.025 0.995 ;
        RECT  5.005 -0.130 5.765 0.130 ;
        RECT  4.745 -0.130 5.005 0.905 ;
        RECT  3.985 -0.130 4.745 0.130 ;
        RECT  3.725 -0.130 3.985 0.905 ;
        RECT  2.965 -0.130 3.725 0.130 ;
        RECT  2.705 -0.130 2.965 0.565 ;
        RECT  0.925 -0.130 2.705 0.130 ;
        RECT  0.665 -0.130 0.925 0.670 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 2.740 6.150 3.000 ;
        RECT  5.765 1.870 6.025 3.000 ;
        RECT  5.005 2.740 5.765 3.000 ;
        RECT  4.745 1.965 5.005 3.000 ;
        RECT  3.985 2.740 4.745 3.000 ;
        RECT  3.725 1.965 3.985 3.000 ;
        RECT  2.965 2.740 3.725 3.000 ;
        RECT  2.705 2.305 2.965 3.000 ;
        RECT  0.925 2.740 2.705 3.000 ;
        RECT  0.665 2.130 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.465 1.355 2.630 1.515 ;
        RECT  1.305 0.385 1.465 2.390 ;
        RECT  1.205 0.385 1.305 1.020 ;
        RECT  1.205 1.760 1.305 2.390 ;
        RECT  0.385 0.860 1.205 1.020 ;
        RECT  0.385 1.760 1.205 1.920 ;
        RECT  0.125 0.395 0.385 1.020 ;
        RECT  0.125 1.760 0.385 2.410 ;
    END
END BUFX16MTH

MACRO BUFX18MTH
    CLASS CORE ;
    FOREIGN BUFX18MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.585 0.425 6.845 2.335 ;
        RECT  5.825 1.050 6.585 1.820 ;
        RECT  5.565 0.425 5.825 2.335 ;
        RECT  4.805 1.050 5.565 1.820 ;
        RECT  4.545 0.425 4.805 2.335 ;
        RECT  3.785 1.050 4.545 1.820 ;
        RECT  3.525 0.420 3.785 2.335 ;
        RECT  3.330 0.745 3.525 2.125 ;
        RECT  2.765 0.745 3.330 1.145 ;
        RECT  2.765 1.735 3.330 2.125 ;
        RECT  2.505 0.420 2.765 1.145 ;
        RECT  2.505 1.735 2.765 2.335 ;
        END
        AntennaDiffArea 2.937 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.375 1.290 1.315 1.580 ;
        END
        AntennaGateArea 0.7592 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 -0.130 6.970 0.130 ;
        RECT  6.075 -0.130 6.335 0.785 ;
        RECT  5.315 -0.130 6.075 0.130 ;
        RECT  5.055 -0.130 5.315 0.785 ;
        RECT  4.295 -0.130 5.055 0.130 ;
        RECT  4.035 -0.130 4.295 0.785 ;
        RECT  3.275 -0.130 4.035 0.130 ;
        RECT  3.015 -0.130 3.275 0.565 ;
        RECT  2.255 -0.130 3.015 0.130 ;
        RECT  1.995 -0.130 2.255 0.955 ;
        RECT  0.385 -0.130 1.995 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 2.740 6.970 3.000 ;
        RECT  6.075 2.095 6.335 3.000 ;
        RECT  5.315 2.740 6.075 3.000 ;
        RECT  5.055 2.095 5.315 3.000 ;
        RECT  4.295 2.740 5.055 3.000 ;
        RECT  4.035 2.095 4.295 3.000 ;
        RECT  3.275 2.740 4.035 3.000 ;
        RECT  3.015 2.305 3.275 3.000 ;
        RECT  2.255 2.740 3.015 3.000 ;
        RECT  1.995 1.775 2.255 3.000 ;
        RECT  0.385 2.740 1.995 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.670 1.355 2.950 1.515 ;
        RECT  1.670 0.420 1.745 1.020 ;
        RECT  1.670 1.790 1.745 2.390 ;
        RECT  1.510 0.420 1.670 2.390 ;
        RECT  1.485 0.420 1.510 1.020 ;
        RECT  1.485 1.790 1.510 2.390 ;
        RECT  0.785 0.860 1.485 1.020 ;
        RECT  0.785 1.790 1.485 1.950 ;
        RECT  0.525 0.605 0.785 1.020 ;
        RECT  0.525 1.790 0.785 2.185 ;
    END
END BUFX18MTH

MACRO BUFX20MTH
    CLASS CORE ;
    FOREIGN BUFX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.485 0.425 6.745 2.335 ;
        RECT  5.815 1.015 6.485 1.855 ;
        RECT  5.555 0.425 5.815 2.335 ;
        RECT  4.795 1.015 5.555 1.855 ;
        RECT  4.535 0.425 4.795 2.335 ;
        RECT  3.775 1.015 4.535 1.855 ;
        RECT  3.515 0.420 3.775 2.335 ;
        RECT  2.585 0.420 3.515 1.020 ;
        RECT  2.585 1.735 3.515 2.335 ;
        END
        AntennaDiffArea 3 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.455 1.290 1.405 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.255 -0.130 7.380 0.130 ;
        RECT  6.995 -0.130 7.255 0.955 ;
        RECT  5.305 -0.130 6.995 0.130 ;
        RECT  5.045 -0.130 5.305 0.665 ;
        RECT  4.285 -0.130 5.045 0.130 ;
        RECT  4.025 -0.130 4.285 0.665 ;
        RECT  2.335 -0.130 4.025 0.130 ;
        RECT  2.075 -0.130 2.335 0.980 ;
        RECT  0.385 -0.130 2.075 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.255 2.740 7.380 3.000 ;
        RECT  6.995 1.915 7.255 3.000 ;
        RECT  5.305 2.740 6.995 3.000 ;
        RECT  5.045 2.165 5.305 3.000 ;
        RECT  4.285 2.740 5.045 3.000 ;
        RECT  4.025 2.165 4.285 3.000 ;
        RECT  2.335 2.740 4.025 3.000 ;
        RECT  2.075 1.795 2.335 3.000 ;
        RECT  0.385 2.740 2.075 3.000 ;
        RECT  0.125 1.795 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.825 1.345 3.095 1.505 ;
        RECT  1.665 0.420 1.825 2.405 ;
        RECT  1.565 0.420 1.665 1.020 ;
        RECT  1.565 1.805 1.665 2.405 ;
        RECT  0.895 0.860 1.565 1.020 ;
        RECT  0.895 1.805 1.565 1.965 ;
        RECT  0.635 0.400 0.895 1.020 ;
        RECT  0.635 1.805 0.895 2.405 ;
    END
END BUFX20MTH

MACRO BUFX24MTH
    CLASS CORE ;
    FOREIGN BUFX24MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.105 0.400 8.365 2.355 ;
        RECT  7.345 1.015 8.105 1.855 ;
        RECT  7.085 0.400 7.345 2.355 ;
        RECT  6.325 1.015 7.085 1.855 ;
        RECT  6.065 0.400 6.325 2.355 ;
        RECT  5.395 1.015 6.065 1.855 ;
        RECT  5.135 0.400 5.395 2.355 ;
        RECT  4.375 1.015 5.135 1.855 ;
        RECT  4.115 0.400 4.375 2.355 ;
        RECT  3.185 0.400 4.115 1.000 ;
        RECT  3.185 1.755 4.115 2.355 ;
        END
        AntennaDiffArea 3.516 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.245 2.085 1.505 ;
        RECT  0.920 1.245 1.130 1.580 ;
        RECT  0.465 1.245 0.920 1.505 ;
        END
        AntennaGateArea 1.001 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.885 -0.130 9.020 0.130 ;
        RECT  8.625 -0.130 8.885 0.975 ;
        RECT  7.855 -0.130 8.625 0.130 ;
        RECT  7.595 -0.130 7.855 0.795 ;
        RECT  6.835 -0.130 7.595 0.130 ;
        RECT  6.575 -0.130 6.835 0.790 ;
        RECT  4.885 -0.130 6.575 0.130 ;
        RECT  4.625 -0.130 4.885 0.795 ;
        RECT  2.935 -0.130 4.625 0.130 ;
        RECT  2.675 -0.130 2.935 1.020 ;
        RECT  1.915 -0.130 2.675 0.130 ;
        RECT  1.655 -0.130 1.915 0.710 ;
        RECT  0.895 -0.130 1.655 0.130 ;
        RECT  0.635 -0.130 0.895 0.710 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.885 2.740 9.020 3.000 ;
        RECT  8.625 1.815 8.885 3.000 ;
        RECT  7.855 2.740 8.625 3.000 ;
        RECT  7.595 2.075 7.855 3.000 ;
        RECT  6.835 2.740 7.595 3.000 ;
        RECT  6.575 2.075 6.835 3.000 ;
        RECT  4.885 2.740 6.575 3.000 ;
        RECT  4.625 2.075 4.885 3.000 ;
        RECT  2.935 2.740 4.625 3.000 ;
        RECT  2.675 1.815 2.935 3.000 ;
        RECT  1.915 2.740 2.675 3.000 ;
        RECT  1.655 2.145 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.145 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.425 1.250 3.765 1.510 ;
        RECT  2.265 0.420 2.425 2.385 ;
        RECT  2.165 0.420 2.265 1.055 ;
        RECT  2.165 1.765 2.265 2.385 ;
        RECT  1.405 0.895 2.165 1.055 ;
        RECT  1.405 1.765 2.165 1.925 ;
        RECT  1.145 0.420 1.405 1.055 ;
        RECT  1.145 1.765 1.405 2.365 ;
        RECT  0.385 0.895 1.145 1.055 ;
        RECT  0.385 1.765 1.145 1.925 ;
        RECT  0.125 0.425 0.385 1.055 ;
        RECT  0.125 1.765 0.385 2.365 ;
    END
END BUFX24MTH

MACRO BUFX2MTH
    CLASS CORE ;
    FOREIGN BUFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.495 0.405 1.540 1.990 ;
        RECT  1.380 0.405 1.495 2.395 ;
        RECT  1.285 0.405 1.380 1.005 ;
        RECT  1.235 1.700 1.380 2.395 ;
        END
        AntennaDiffArea 0.524 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 1.185 0.760 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 -0.130 1.640 0.130 ;
        RECT  0.695 -0.130 0.955 0.645 ;
        RECT  0.355 -0.130 0.695 0.300 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 2.740 1.640 3.000 ;
        RECT  0.695 1.880 0.955 3.000 ;
        RECT  0.405 2.740 0.695 3.000 ;
        RECT  0.145 2.570 0.405 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.100 1.210 1.200 1.470 ;
        RECT  0.940 0.845 1.100 1.470 ;
        RECT  0.405 0.845 0.940 1.005 ;
        RECT  0.260 0.745 0.405 1.005 ;
        RECT  0.260 1.755 0.355 2.015 ;
        RECT  0.100 0.745 0.260 2.015 ;
    END
END BUFX2MTH

MACRO BUFX32MTH
    CLASS CORE ;
    FOREIGN BUFX32MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.985 0.400 11.245 2.355 ;
        RECT  10.225 1.015 10.985 1.855 ;
        RECT  9.965 0.400 10.225 2.355 ;
        RECT  9.205 1.015 9.965 1.855 ;
        RECT  8.945 0.400 9.205 2.355 ;
        RECT  8.185 1.015 8.945 1.855 ;
        RECT  7.925 0.400 8.185 2.355 ;
        RECT  7.165 1.015 7.925 1.855 ;
        RECT  6.905 0.400 7.165 2.355 ;
        RECT  6.235 1.015 6.905 1.855 ;
        RECT  5.975 0.400 6.235 2.355 ;
        RECT  5.215 1.015 5.975 1.855 ;
        RECT  4.955 0.400 5.215 2.355 ;
        RECT  4.025 0.400 4.955 1.000 ;
        RECT  4.025 1.755 4.955 2.355 ;
        END
        AntennaDiffArea 4.688 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.245 2.755 1.505 ;
        RECT  1.740 1.245 1.950 1.580 ;
        RECT  0.795 1.245 1.740 1.505 ;
        END
        AntennaGateArea 1.4014 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.755 -0.130 11.890 0.130 ;
        RECT  11.495 -0.130 11.755 0.975 ;
        RECT  10.735 -0.130 11.495 0.130 ;
        RECT  10.475 -0.130 10.735 0.795 ;
        RECT  9.715 -0.130 10.475 0.130 ;
        RECT  9.455 -0.130 9.715 0.800 ;
        RECT  8.695 -0.130 9.455 0.130 ;
        RECT  8.435 -0.130 8.695 0.795 ;
        RECT  7.675 -0.130 8.435 0.130 ;
        RECT  7.415 -0.130 7.675 0.790 ;
        RECT  5.725 -0.130 7.415 0.130 ;
        RECT  5.465 -0.130 5.725 0.795 ;
        RECT  3.775 -0.130 5.465 0.130 ;
        RECT  3.515 -0.130 3.775 1.020 ;
        RECT  0.895 -0.130 3.515 0.130 ;
        RECT  0.635 -0.130 0.895 0.710 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.755 2.740 11.890 3.000 ;
        RECT  11.495 1.860 11.755 3.000 ;
        RECT  10.735 2.740 11.495 3.000 ;
        RECT  10.475 2.075 10.735 3.000 ;
        RECT  9.715 2.740 10.475 3.000 ;
        RECT  9.455 2.075 9.715 3.000 ;
        RECT  8.695 2.740 9.455 3.000 ;
        RECT  8.435 2.075 8.695 3.000 ;
        RECT  7.675 2.740 8.435 3.000 ;
        RECT  7.415 2.075 7.675 3.000 ;
        RECT  5.725 2.740 7.415 3.000 ;
        RECT  5.465 2.075 5.725 3.000 ;
        RECT  3.775 2.740 5.465 3.000 ;
        RECT  3.515 1.815 3.775 3.000 ;
        RECT  0.895 2.740 3.515 3.000 ;
        RECT  0.635 2.145 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.835 1.250 4.775 1.510 ;
        RECT  3.265 1.305 3.835 1.465 ;
        RECT  3.105 0.420 3.265 2.385 ;
        RECT  3.005 0.420 3.105 1.050 ;
        RECT  3.005 1.765 3.105 2.385 ;
        RECT  2.335 0.890 3.005 1.050 ;
        RECT  2.335 1.765 3.005 1.925 ;
        RECT  2.075 0.420 2.335 1.050 ;
        RECT  2.075 1.765 2.335 2.365 ;
        RECT  1.405 0.890 2.075 1.050 ;
        RECT  1.405 1.765 2.075 1.925 ;
        RECT  1.145 0.425 1.405 1.050 ;
        RECT  1.145 1.765 1.405 2.365 ;
        RECT  0.385 0.890 1.145 1.050 ;
        RECT  0.385 1.765 1.145 1.925 ;
        RECT  0.125 0.420 0.385 1.050 ;
        RECT  0.125 1.765 0.385 2.365 ;
    END
END BUFX32MTH

MACRO BUFX3MTH
    CLASS CORE ;
    FOREIGN BUFX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 1.290 1.950 1.580 ;
        RECT  1.610 0.875 1.770 1.935 ;
        RECT  1.405 0.875 1.610 1.035 ;
        RECT  1.405 1.775 1.610 1.935 ;
        RECT  1.145 0.575 1.405 1.035 ;
        RECT  1.145 1.775 1.405 2.105 ;
        END
        AntennaDiffArea 0.472 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 0.880 0.915 1.255 ;
        END
        AntennaGateArea 0.1326 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 -0.130 2.050 0.130 ;
        RECT  1.655 -0.130 1.915 0.695 ;
        RECT  0.895 -0.130 1.655 0.130 ;
        RECT  0.635 -0.130 0.895 0.700 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 2.740 2.050 3.000 ;
        RECT  1.655 2.115 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.605 1.955 0.895 3.000 ;
        RECT  0.265 2.570 0.605 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.110 1.235 1.370 1.595 ;
        RECT  0.385 1.435 1.110 1.595 ;
        RECT  0.285 0.455 0.385 0.715 ;
        RECT  0.285 1.435 0.385 2.055 ;
        RECT  0.125 0.455 0.285 2.055 ;
    END
END BUFX3MTH

MACRO BUFX4MTH
    CLASS CORE ;
    FOREIGN BUFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 0.810 1.550 1.990 ;
        RECT  1.370 0.380 1.405 2.400 ;
        RECT  1.145 0.380 1.370 0.990 ;
        RECT  1.145 1.690 1.370 2.400 ;
        END
        AntennaDiffArea 0.586 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.260 0.555 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 -0.130 2.050 0.130 ;
        RECT  1.655 -0.130 1.915 0.640 ;
        RECT  0.895 -0.130 1.655 0.130 ;
        RECT  0.635 -0.130 0.895 0.735 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 2.740 2.050 3.000 ;
        RECT  1.655 2.170 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.125 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.905 1.250 1.185 1.510 ;
        RECT  0.745 0.915 0.905 1.920 ;
        RECT  0.385 0.915 0.745 1.075 ;
        RECT  0.385 1.760 0.745 1.920 ;
        RECT  0.125 0.765 0.385 1.075 ;
        RECT  0.125 1.760 0.385 2.380 ;
    END
END BUFX4MTH

MACRO BUFX5MTH
    CLASS CORE ;
    FOREIGN BUFX5MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.285 0.715 2.335 0.975 ;
        RECT  2.285 1.685 2.335 1.945 ;
        RECT  2.075 0.715 2.285 1.945 ;
        RECT  1.540 1.265 2.075 1.475 ;
        RECT  1.385 0.820 1.540 1.995 ;
        RECT  1.330 0.400 1.385 2.415 ;
        RECT  1.125 0.400 1.330 1.000 ;
        RECT  1.125 1.815 1.330 2.415 ;
        END
        AntennaDiffArea 0.885 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.255 0.555 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 -0.130 2.460 0.130 ;
        RECT  1.665 -0.130 2.265 0.300 ;
        RECT  0.000 -0.130 1.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 2.740 2.460 3.000 ;
        RECT  1.665 2.570 2.265 3.000 ;
        RECT  0.000 2.740 1.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.945 1.205 1.150 1.465 ;
        RECT  0.785 0.835 0.945 1.920 ;
        RECT  0.385 0.835 0.785 0.995 ;
        RECT  0.385 1.760 0.785 1.920 ;
        RECT  0.125 0.395 0.385 0.995 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END BUFX5MTH

MACRO BUFX6MTH
    CLASS CORE ;
    FOREIGN BUFX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.475 0.405 2.745 1.035 ;
        RECT  2.475 1.615 2.745 2.305 ;
        RECT  2.395 0.765 2.475 1.035 ;
        RECT  2.395 1.615 2.475 1.885 ;
        RECT  2.115 0.765 2.395 1.885 ;
        RECT  1.735 0.765 2.115 1.035 ;
        RECT  1.735 1.615 2.115 1.885 ;
        RECT  1.465 0.380 1.735 1.035 ;
        RECT  1.465 1.615 1.735 2.400 ;
        END
        AntennaDiffArea 1.11 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.210 0.905 1.470 ;
        RECT  0.100 1.210 0.310 1.580 ;
        END
        AntennaGateArea 0.26 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 -0.130 2.870 0.130 ;
        RECT  1.975 -0.130 2.235 0.585 ;
        RECT  1.110 -0.130 1.975 0.130 ;
        RECT  0.170 -0.130 1.110 0.300 ;
        RECT  0.000 -0.130 0.170 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 2.740 2.870 3.000 ;
        RECT  1.975 2.065 2.235 3.000 ;
        RECT  1.100 2.740 1.975 3.000 ;
        RECT  0.160 2.570 1.100 3.000 ;
        RECT  0.000 2.740 0.160 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.285 1.215 1.895 1.435 ;
        RECT  1.125 0.850 1.285 1.940 ;
        RECT  0.785 0.850 1.125 1.010 ;
        RECT  0.785 1.780 1.125 1.940 ;
        RECT  0.525 0.750 0.785 1.010 ;
        RECT  0.525 1.780 0.785 2.040 ;
    END
END BUFX6MTH

MACRO BUFX8MTH
    CLASS CORE ;
    FOREIGN BUFX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.445 0.670 2.785 1.110 ;
        RECT  2.445 1.730 2.785 2.170 ;
        RECT  2.380 0.770 2.445 1.110 ;
        RECT  2.380 1.730 2.445 2.070 ;
        RECT  1.930 0.770 2.380 2.070 ;
        RECT  1.765 0.770 1.930 1.110 ;
        RECT  1.760 1.730 1.930 2.070 ;
        RECT  1.425 0.380 1.765 1.110 ;
        RECT  1.420 1.730 1.760 2.400 ;
        END
        AntennaDiffArea 1.131 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.245 0.875 1.505 ;
        RECT  0.275 1.245 0.720 1.580 ;
        END
        AntennaGateArea 0.3445 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 -0.130 3.280 0.130 ;
        RECT  2.895 -0.130 3.155 0.300 ;
        RECT  2.235 -0.130 2.895 0.130 ;
        RECT  1.975 -0.130 2.235 0.565 ;
        RECT  0.385 -0.130 1.975 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.895 2.570 3.155 3.000 ;
        RECT  2.235 2.740 2.895 3.000 ;
        RECT  1.975 2.280 2.235 3.000 ;
        RECT  0.385 2.740 1.975 3.000 ;
        RECT  0.125 2.535 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.215 1.290 1.655 1.550 ;
        RECT  1.055 0.905 1.215 1.930 ;
        RECT  0.795 0.905 1.055 1.065 ;
        RECT  0.795 1.770 1.055 1.930 ;
        RECT  0.635 0.630 0.795 1.065 ;
        RECT  0.535 1.770 0.795 2.140 ;
        RECT  0.535 0.630 0.635 0.890 ;
    END
END BUFX8MTH

MACRO CLKAND2X12MTH
    CLASS CORE ;
    FOREIGN CLKAND2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.025 1.805 5.105 2.405 ;
        RECT  5.025 0.465 5.080 1.005 ;
        RECT  4.405 0.465 5.025 2.405 ;
        RECT  3.680 0.465 4.405 1.005 ;
        RECT  2.960 1.805 4.405 2.405 ;
        END
        AntennaDiffArea 1.461 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.070 2.410 1.745 ;
        RECT  1.110 1.585 2.110 1.745 ;
        RECT  0.950 1.065 1.110 1.745 ;
        RECT  0.865 1.065 0.950 1.325 ;
        END
        AntennaGateArea 0.3666 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 0.920 1.760 1.250 ;
        END
        AntennaGateArea 0.3666 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.515 -0.130 5.740 0.130 ;
        RECT  4.255 -0.130 4.515 0.250 ;
        RECT  3.380 -0.130 4.255 0.130 ;
        RECT  3.120 -0.130 3.380 0.840 ;
        RECT  2.440 -0.130 3.120 0.300 ;
        RECT  0.960 -0.130 2.440 0.130 ;
        RECT  0.700 -0.130 0.960 0.790 ;
        RECT  0.000 -0.130 0.700 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 1.885 5.615 3.000 ;
        RECT  0.760 2.740 5.355 3.000 ;
        RECT  0.500 1.940 0.760 3.000 ;
        RECT  0.000 2.740 0.500 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.750 1.225 4.020 1.485 ;
        RECT  2.590 0.580 2.750 2.095 ;
        RECT  1.550 0.580 2.590 0.740 ;
        RECT  2.230 1.935 2.590 2.095 ;
        RECT  1.970 1.935 2.230 2.435 ;
        RECT  1.300 1.935 1.970 2.095 ;
        RECT  1.040 1.935 1.300 2.435 ;
    END
END CLKAND2X12MTH

MACRO CLKAND2X16MTH
    CLASS CORE ;
    FOREIGN CLKAND2X16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.585 1.085 6.845 2.325 ;
        RECT  5.825 1.085 6.585 1.785 ;
        RECT  5.565 1.085 5.825 2.325 ;
        RECT  4.800 1.085 5.565 1.785 ;
        RECT  4.540 1.085 4.800 2.325 ;
        RECT  4.265 1.085 4.540 1.785 ;
        RECT  4.265 0.415 4.505 0.675 ;
        RECT  3.775 0.415 4.265 1.785 ;
        RECT  3.565 0.415 3.775 2.325 ;
        RECT  3.315 0.415 3.565 0.675 ;
        RECT  3.515 1.725 3.565 2.325 ;
        END
        AntennaDiffArea 1.956 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.795 1.195 2.895 1.455 ;
        RECT  2.635 1.195 2.795 1.745 ;
        RECT  1.225 1.585 2.635 1.745 ;
        RECT  0.920 1.205 1.225 1.745 ;
        END
        AntennaGateArea 0.5174 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.245 2.305 1.405 ;
        RECT  1.705 0.865 1.950 1.405 ;
        RECT  0.675 0.865 1.705 1.025 ;
        RECT  0.515 0.865 0.675 1.495 ;
        END
        AntennaGateArea 0.5174 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.015 -0.130 6.970 0.130 ;
        RECT  4.755 -0.130 5.015 0.755 ;
        RECT  3.065 -0.130 4.755 0.130 ;
        RECT  2.805 -0.130 3.065 0.665 ;
        RECT  1.285 -0.130 2.805 0.130 ;
        RECT  1.025 -0.130 1.285 0.640 ;
        RECT  0.000 -0.130 1.025 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 2.740 6.970 3.000 ;
        RECT  6.075 1.965 6.335 3.000 ;
        RECT  5.310 2.740 6.075 3.000 ;
        RECT  5.050 1.965 5.310 3.000 ;
        RECT  4.290 2.740 5.050 3.000 ;
        RECT  4.030 1.965 4.290 3.000 ;
        RECT  3.265 2.740 4.030 3.000 ;
        RECT  3.005 2.275 3.265 3.000 ;
        RECT  0.385 2.740 3.005 3.000 ;
        RECT  0.125 1.905 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.240 1.115 3.385 1.375 ;
        RECT  3.080 0.855 3.240 2.090 ;
        RECT  2.290 0.855 3.080 1.015 ;
        RECT  2.755 1.930 3.080 2.090 ;
        RECT  2.495 1.930 2.755 2.465 ;
        RECT  1.825 1.930 2.495 2.090 ;
        RECT  2.130 0.420 2.290 1.015 ;
        RECT  1.925 0.420 2.130 0.680 ;
        RECT  1.565 1.930 1.825 2.465 ;
        RECT  0.895 1.930 1.565 2.090 ;
        RECT  0.635 1.930 0.895 2.465 ;
    END
END CLKAND2X16MTH

MACRO CLKAND2X2MTH
    CLASS CORE ;
    FOREIGN CLKAND2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 1.290 1.950 1.580 ;
        RECT  1.715 0.665 1.875 2.345 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 0.920 1.170 1.500 ;
        END
        AntennaGateArea 0.0689 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.280 0.470 1.635 ;
        END
        AntennaGateArea 0.0689 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 -0.130 2.050 0.130 ;
        RECT  1.245 -0.130 1.845 0.300 ;
        RECT  1.065 -0.130 1.245 0.130 ;
        RECT  0.125 -0.130 1.065 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 2.740 2.050 3.000 ;
        RECT  0.260 2.290 1.200 3.000 ;
        RECT  0.000 2.740 0.260 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.375 0.580 1.535 1.895 ;
        RECT  0.385 0.580 1.375 0.740 ;
        RECT  0.955 1.735 1.375 1.895 ;
        RECT  0.685 1.735 0.955 1.995 ;
        RECT  0.175 0.580 0.385 0.875 ;
        RECT  0.125 0.615 0.175 0.875 ;
    END
END CLKAND2X2MTH

MACRO CLKAND2X3MTH
    CLASS CORE ;
    FOREIGN CLKAND2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.870 0.705 2.030 1.990 ;
        RECT  1.745 0.705 1.870 0.965 ;
        RECT  1.650 1.700 1.870 2.310 ;
        END
        AntennaDiffArea 0.435 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.845 1.190 1.130 1.725 ;
        END
        AntennaGateArea 0.0962 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.245 0.640 1.580 ;
        END
        AntennaGateArea 0.0962 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 -0.130 2.460 0.130 ;
        RECT  1.915 -0.130 2.175 0.300 ;
        RECT  1.465 -0.130 1.915 0.130 ;
        RECT  0.865 -0.130 1.465 0.300 ;
        RECT  0.575 -0.130 0.865 0.130 ;
        RECT  0.315 -0.130 0.575 0.300 ;
        RECT  0.000 -0.130 0.315 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 2.740 2.460 3.000 ;
        RECT  2.060 2.570 2.320 3.000 ;
        RECT  1.310 2.740 2.060 3.000 ;
        RECT  0.710 2.570 1.310 3.000 ;
        RECT  0.385 2.740 0.710 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.470 1.225 1.690 1.485 ;
        RECT  1.310 0.810 1.470 2.070 ;
        RECT  0.500 0.810 1.310 0.970 ;
        RECT  0.860 1.910 1.310 2.070 ;
        RECT  0.600 1.910 0.860 2.170 ;
        RECT  0.240 0.710 0.500 0.970 ;
    END
END CLKAND2X3MTH

MACRO CLKAND2X4MTH
    CLASS CORE ;
    FOREIGN CLKAND2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 0.460 1.950 1.795 ;
        RECT  1.740 0.460 1.840 2.365 ;
        RECT  1.565 0.460 1.740 0.720 ;
        RECT  1.660 1.615 1.740 2.365 ;
        RECT  1.565 2.105 1.660 2.365 ;
        END
        AntennaDiffArea 0.541 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.740 1.240 1.130 1.580 ;
        END
        AntennaGateArea 0.13 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 1.240 0.555 1.500 ;
        RECT  0.100 1.240 0.355 1.990 ;
        END
        AntennaGateArea 0.13 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 -0.130 2.460 0.130 ;
        RECT  2.070 -0.130 2.330 0.300 ;
        RECT  1.260 -0.130 2.070 0.130 ;
        RECT  1.000 -0.130 1.260 0.665 ;
        RECT  0.320 -0.130 1.000 0.300 ;
        RECT  0.000 -0.130 0.320 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  2.075 1.965 2.335 3.000 ;
        RECT  1.315 2.740 2.075 3.000 ;
        RECT  1.055 2.105 1.315 3.000 ;
        RECT  0.000 2.740 1.055 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.480 1.170 1.550 1.430 ;
        RECT  1.320 0.900 1.480 1.920 ;
        RECT  0.385 0.900 1.320 1.060 ;
        RECT  0.800 1.760 1.320 1.920 ;
        RECT  0.540 1.760 0.800 2.260 ;
        RECT  0.125 0.755 0.385 1.060 ;
    END
END CLKAND2X4MTH

MACRO CLKAND2X6MTH
    CLASS CORE ;
    FOREIGN CLKAND2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 0.810 2.775 1.990 ;
        RECT  2.505 0.590 2.550 2.365 ;
        RECT  2.280 0.590 2.505 1.080 ;
        RECT  2.280 1.700 2.505 2.365 ;
        RECT  0.335 2.105 2.280 2.365 ;
        RECT  0.135 1.765 0.335 2.365 ;
        END
        AntennaDiffArea 0.798 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.880 1.620 1.580 ;
        END
        AntennaGateArea 0.1911 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 0.880 1.150 1.585 ;
        END
        AntennaGateArea 0.1911 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 -0.130 3.280 0.130 ;
        RECT  2.825 -0.130 3.085 0.630 ;
        RECT  1.905 -0.130 2.825 0.130 ;
        RECT  1.645 -0.130 1.905 0.300 ;
        RECT  0.445 -0.130 1.645 0.130 ;
        RECT  0.185 -0.130 0.445 0.300 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.085 2.740 3.280 3.000 ;
        RECT  2.825 2.230 3.085 3.000 ;
        RECT  2.005 2.740 2.825 3.000 ;
        RECT  1.745 2.570 2.005 3.000 ;
        RECT  0.925 2.740 1.745 3.000 ;
        RECT  0.665 2.570 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.965 1.260 2.325 1.520 ;
        RECT  1.805 0.540 1.965 1.925 ;
        RECT  0.695 0.540 1.805 0.700 ;
        RECT  0.675 1.765 1.805 1.925 ;
        RECT  0.515 1.365 0.675 1.925 ;
        RECT  0.295 1.365 0.515 1.525 ;
    END
END CLKAND2X6MTH

MACRO CLKAND2X8MTH
    CLASS CORE ;
    FOREIGN CLKAND2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.730 1.720 3.915 2.440 ;
        RECT  3.565 0.625 3.730 2.440 ;
        RECT  3.380 0.625 3.565 2.070 ;
        RECT  2.545 0.625 3.380 0.975 ;
        RECT  2.895 1.720 3.380 2.070 ;
        RECT  2.545 1.720 2.895 2.405 ;
        END
        AntennaDiffArea 0.92 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.705 1.240 1.970 1.745 ;
        RECT  0.725 1.585 1.705 1.745 ;
        RECT  0.565 1.245 0.725 1.745 ;
        RECT  0.465 1.245 0.565 1.505 ;
        END
        AntennaGateArea 0.2587 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.355 1.405 ;
        END
        AntennaGateArea 0.2587 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.510 0.130 ;
        RECT  3.035 -0.130 3.975 0.300 ;
        RECT  2.165 -0.130 3.035 0.130 ;
        RECT  1.905 -0.130 2.165 0.250 ;
        RECT  0.805 -0.130 1.905 0.130 ;
        RECT  0.205 -0.130 0.805 0.300 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.965 4.385 3.000 ;
        RECT  3.360 2.740 4.125 3.000 ;
        RECT  3.100 2.255 3.360 3.000 ;
        RECT  2.335 2.740 3.100 3.000 ;
        RECT  2.075 2.275 2.335 3.000 ;
        RECT  0.385 2.740 2.075 3.000 ;
        RECT  0.125 1.935 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.345 1.225 3.190 1.485 ;
        RECT  2.185 0.525 2.345 2.095 ;
        RECT  1.055 0.525 2.185 0.685 ;
        RECT  1.825 1.935 2.185 2.095 ;
        RECT  1.565 1.935 1.825 2.435 ;
        RECT  0.895 1.935 1.565 2.095 ;
        RECT  0.635 1.935 0.895 2.435 ;
    END
END CLKAND2X8MTH

MACRO CLKBUFX12MTH
    CLASS CORE ;
    FOREIGN CLKBUFX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 1.735 3.875 2.335 ;
        RECT  3.105 1.735 3.615 2.115 ;
        RECT  2.945 0.765 3.105 2.115 ;
        RECT  2.845 0.765 2.945 2.335 ;
        RECT  2.685 0.770 2.845 2.335 ;
        RECT  2.355 0.770 2.685 2.115 ;
        RECT  1.990 0.770 2.355 1.150 ;
        RECT  1.925 1.735 2.355 2.115 ;
        RECT  1.730 0.425 1.990 1.150 ;
        RECT  1.665 1.735 1.925 2.335 ;
        END
        AntennaDiffArea 1.41 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.250 0.585 1.580 ;
        END
        AntennaGateArea 0.2899 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 -0.130 4.510 0.130 ;
        RECT  3.415 -0.130 4.015 1.025 ;
        RECT  3.105 -0.130 3.415 0.130 ;
        RECT  2.845 -0.130 3.105 0.385 ;
        RECT  2.560 -0.130 2.845 0.130 ;
        RECT  2.300 -0.130 2.560 0.590 ;
        RECT  1.420 -0.130 2.300 0.130 ;
        RECT  1.160 -0.130 1.420 1.025 ;
        RECT  0.725 -0.130 1.160 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.890 4.385 3.000 ;
        RECT  2.435 2.740 4.125 3.000 ;
        RECT  2.175 2.305 2.435 3.000 ;
        RECT  1.410 2.740 2.175 3.000 ;
        RECT  1.150 1.825 1.410 3.000 ;
        RECT  0.385 2.740 1.150 3.000 ;
        RECT  0.125 1.825 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.935 1.355 2.095 1.515 ;
        RECT  0.775 0.765 0.935 2.425 ;
        RECT  0.610 0.765 0.775 1.025 ;
        RECT  0.635 1.825 0.775 2.425 ;
    END
END CLKBUFX12MTH

MACRO CLKBUFX16MTH
    CLASS CORE ;
    FOREIGN CLKBUFX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 1.385 5.205 2.355 ;
        RECT  4.245 1.385 4.945 1.785 ;
        RECT  3.385 0.465 4.445 0.865 ;
        RECT  3.985 1.385 4.245 2.335 ;
        RECT  3.385 1.385 3.985 1.785 ;
        RECT  3.305 0.465 3.385 1.785 ;
        RECT  3.045 0.465 3.305 2.335 ;
        RECT  2.765 0.465 3.045 1.785 ;
        RECT  1.995 0.465 2.765 0.865 ;
        RECT  2.285 1.385 2.765 1.785 ;
        RECT  2.025 1.385 2.285 2.335 ;
        END
        AntennaDiffArea 1.956 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.325 1.290 0.865 1.580 ;
        END
        AntennaGateArea 0.3913 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.025 -0.130 5.330 0.130 ;
        RECT  4.765 -0.130 5.025 0.825 ;
        RECT  4.555 -0.130 4.765 0.130 ;
        RECT  3.615 -0.130 4.555 0.250 ;
        RECT  2.795 -0.130 3.615 0.130 ;
        RECT  2.535 -0.130 2.795 0.250 ;
        RECT  1.715 -0.130 2.535 0.130 ;
        RECT  1.455 -0.130 1.715 0.640 ;
        RECT  0.635 -0.130 1.455 0.130 ;
        RECT  0.375 -0.130 0.635 0.825 ;
        RECT  0.000 -0.130 0.375 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.795 2.740 5.330 3.000 ;
        RECT  2.535 1.965 2.795 3.000 ;
        RECT  0.785 2.740 2.535 3.000 ;
        RECT  0.185 2.485 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.325 1.045 2.430 1.205 ;
        RECT  1.175 0.860 1.325 2.390 ;
        RECT  1.165 0.530 1.175 2.390 ;
        RECT  0.915 0.530 1.165 1.020 ;
        RECT  1.065 1.760 1.165 2.390 ;
        RECT  0.385 1.760 1.065 1.920 ;
        RECT  0.125 1.760 0.385 2.020 ;
    END
END CLKBUFX16MTH

MACRO CLKBUFX1MTH
    CLASS CORE ;
    FOREIGN CLKBUFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.765 1.540 2.050 ;
        RECT  1.255 0.765 1.330 1.025 ;
        RECT  1.240 1.770 1.330 2.050 ;
        END
        AntennaDiffArea 0.281 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.585 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 -0.130 1.640 0.130 ;
        RECT  0.335 -0.130 1.275 0.510 ;
        RECT  0.000 -0.130 0.335 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.495 2.740 1.640 3.000 ;
        RECT  1.235 2.485 1.495 3.000 ;
        RECT  0.955 2.740 1.235 3.000 ;
        RECT  0.695 2.195 0.955 3.000 ;
        RECT  0.405 2.740 0.695 3.000 ;
        RECT  0.145 2.485 0.405 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.060 1.240 1.150 1.500 ;
        RECT  0.900 0.950 1.060 1.920 ;
        RECT  0.385 0.950 0.900 1.110 ;
        RECT  0.415 1.760 0.900 1.920 ;
        RECT  0.155 1.760 0.415 2.085 ;
        RECT  0.125 0.765 0.385 1.110 ;
    END
END CLKBUFX1MTH

MACRO CLKBUFX20MTH
    CLASS CORE ;
    FOREIGN CLKBUFX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.600 0.425 5.920 2.495 ;
        RECT  4.925 0.835 5.600 1.675 ;
        RECT  4.665 0.430 4.925 2.460 ;
        RECT  3.845 0.430 4.665 2.010 ;
        RECT  3.585 0.430 3.845 2.460 ;
        RECT  3.540 0.430 3.585 2.010 ;
        RECT  2.375 0.430 3.540 0.910 ;
        RECT  2.810 1.510 3.540 2.010 ;
        RECT  2.550 1.510 2.810 2.460 ;
        END
        AntennaDiffArea 2.276 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.415 1.160 1.155 1.410 ;
        RECT  0.100 1.160 0.415 1.580 ;
        END
        AntennaGateArea 0.4849 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.640 ;
        RECT  5.355 -0.130 6.175 0.130 ;
        RECT  5.095 -0.130 5.355 0.250 ;
        RECT  4.275 -0.130 5.095 0.130 ;
        RECT  4.015 -0.130 4.275 0.250 ;
        RECT  2.135 -0.130 4.015 0.130 ;
        RECT  1.875 -0.130 2.135 0.640 ;
        RECT  1.035 -0.130 1.875 0.130 ;
        RECT  0.775 -0.130 1.035 0.640 ;
        RECT  0.000 -0.130 0.775 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.885 6.435 3.000 ;
        RECT  4.385 2.740 6.175 3.000 ;
        RECT  4.125 2.230 4.385 3.000 ;
        RECT  2.270 2.740 4.125 3.000 ;
        RECT  1.330 2.490 2.270 3.000 ;
        RECT  0.385 2.740 1.330 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.870 1.090 3.205 1.330 ;
        RECT  1.610 1.090 1.870 2.165 ;
        RECT  1.575 1.090 1.610 1.800 ;
        RECT  1.375 0.505 1.575 1.800 ;
        RECT  1.315 0.505 1.375 0.980 ;
        RECT  0.925 1.600 1.375 1.800 ;
        RECT  0.495 0.820 1.315 0.980 ;
        RECT  0.665 1.600 0.925 2.335 ;
        RECT  0.335 0.515 0.495 0.980 ;
        RECT  0.235 0.515 0.335 0.775 ;
    END
END CLKBUFX20MTH

MACRO CLKBUFX24MTH
    CLASS CORE ;
    FOREIGN CLKBUFX24MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.910 1.565 6.410 2.165 ;
        RECT  4.815 0.435 5.910 2.165 ;
        RECT  2.405 0.435 4.815 0.915 ;
        RECT  2.405 1.565 4.815 2.165 ;
        END
        AntennaDiffArea 2.728 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 1.115 1.295 1.375 ;
        RECT  0.355 1.115 0.955 1.580 ;
        END
        AntennaGateArea 0.5837 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.790 -0.130 6.970 0.130 ;
        RECT  6.190 -0.130 6.790 0.725 ;
        RECT  5.370 -0.130 6.190 0.130 ;
        RECT  5.110 -0.130 5.370 0.250 ;
        RECT  4.290 -0.130 5.110 0.130 ;
        RECT  4.030 -0.130 4.290 0.250 ;
        RECT  3.210 -0.130 4.030 0.130 ;
        RECT  2.950 -0.130 3.210 0.250 ;
        RECT  2.125 -0.130 2.950 0.130 ;
        RECT  1.865 -0.130 2.125 0.590 ;
        RECT  1.045 -0.130 1.865 0.130 ;
        RECT  0.785 -0.130 1.045 0.590 ;
        RECT  0.000 -0.130 0.785 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 2.570 6.845 3.000 ;
        RECT  1.130 2.740 6.585 3.000 ;
        RECT  0.190 2.570 1.130 3.000 ;
        RECT  0.000 2.740 0.190 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.725 1.135 4.535 1.295 ;
        RECT  1.585 0.770 1.725 2.360 ;
        RECT  1.565 0.485 1.585 2.360 ;
        RECT  1.325 0.485 1.565 0.930 ;
        RECT  1.465 1.760 1.565 2.360 ;
        RECT  0.785 1.760 1.465 1.920 ;
        RECT  0.505 0.770 1.325 0.930 ;
        RECT  0.525 1.760 0.785 2.090 ;
        RECT  0.245 0.485 0.505 0.930 ;
    END
END CLKBUFX24MTH

MACRO CLKBUFX2MTH
    CLASS CORE ;
    FOREIGN CLKBUFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.360 0.570 1.540 2.290 ;
        RECT  1.255 0.570 1.360 0.830 ;
        RECT  1.255 1.690 1.360 2.290 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.585 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.960 -0.130 1.640 0.130 ;
        RECT  0.700 -0.130 0.960 0.770 ;
        RECT  0.355 -0.130 0.700 0.320 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.970 2.740 1.640 3.000 ;
        RECT  0.710 2.145 0.970 3.000 ;
        RECT  0.370 2.445 0.710 3.000 ;
        RECT  0.000 2.740 0.370 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.060 1.170 1.125 1.430 ;
        RECT  0.900 0.950 1.060 1.920 ;
        RECT  0.385 0.950 0.900 1.110 ;
        RECT  0.420 1.760 0.900 1.920 ;
        RECT  0.160 1.760 0.420 2.020 ;
        RECT  0.225 0.570 0.385 1.110 ;
        RECT  0.125 0.570 0.225 0.830 ;
    END
END CLKBUFX2MTH

MACRO CLKBUFX32MTH
    CLASS CORE ;
    FOREIGN CLKBUFX32MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.785 0.425 8.075 1.760 ;
        RECT  7.625 0.860 7.785 1.760 ;
        RECT  7.245 0.860 7.625 2.370 ;
        RECT  7.025 0.860 7.245 1.940 ;
        RECT  6.705 0.490 7.025 1.940 ;
        RECT  6.635 0.860 6.705 1.940 ;
        RECT  6.375 0.860 6.635 2.485 ;
        RECT  6.005 0.860 6.375 1.940 ;
        RECT  5.705 0.490 6.005 1.940 ;
        RECT  5.685 0.490 5.705 2.485 ;
        RECT  5.445 0.860 5.685 2.485 ;
        RECT  4.985 0.860 5.445 1.940 ;
        RECT  4.775 0.480 4.985 1.940 ;
        RECT  4.665 0.480 4.775 2.485 ;
        RECT  4.515 0.860 4.665 2.485 ;
        RECT  3.975 0.860 4.515 1.940 ;
        RECT  3.695 0.480 3.975 1.940 ;
        RECT  3.470 0.480 3.695 2.485 ;
        RECT  2.595 0.480 3.470 0.890 ;
        RECT  3.435 1.410 3.470 2.485 ;
        RECT  2.765 1.410 3.435 1.940 ;
        RECT  2.505 1.410 2.765 2.485 ;
        END
        AntennaDiffArea 3.574 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 1.045 1.415 1.305 ;
        RECT  0.475 1.045 0.735 1.580 ;
        END
        AntennaGateArea 0.7605 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 -0.130 8.200 0.130 ;
        RECT  7.275 -0.130 7.535 0.680 ;
        RECT  6.485 -0.130 7.275 0.130 ;
        RECT  6.225 -0.130 6.485 0.635 ;
        RECT  5.465 -0.130 6.225 0.130 ;
        RECT  5.205 -0.130 5.465 0.635 ;
        RECT  4.445 -0.130 5.205 0.130 ;
        RECT  4.185 -0.130 4.445 0.635 ;
        RECT  3.395 -0.130 4.185 0.130 ;
        RECT  3.135 -0.130 3.395 0.300 ;
        RECT  2.345 -0.130 3.135 0.130 ;
        RECT  2.085 -0.130 2.345 0.670 ;
        RECT  0.395 -0.130 2.085 0.130 ;
        RECT  0.135 -0.130 0.395 0.665 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 2.740 8.200 3.000 ;
        RECT  7.815 1.965 8.075 3.000 ;
        RECT  4.235 2.740 7.815 3.000 ;
        RECT  3.975 2.140 4.235 3.000 ;
        RECT  0.395 2.740 3.975 3.000 ;
        RECT  0.135 1.915 0.395 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.755 1.070 3.275 1.230 ;
        RECT  1.755 0.435 1.835 0.695 ;
        RECT  1.755 1.715 1.835 2.315 ;
        RECT  1.595 0.435 1.755 2.315 ;
        RECT  1.575 0.435 1.595 0.715 ;
        RECT  1.575 1.715 1.595 2.315 ;
        RECT  0.905 0.555 1.575 0.715 ;
        RECT  0.905 1.780 1.575 1.940 ;
        RECT  0.645 0.455 0.905 0.715 ;
        RECT  0.645 1.780 0.905 2.380 ;
    END
END CLKBUFX32MTH

MACRO CLKBUFX3MTH
    CLASS CORE ;
    FOREIGN CLKBUFX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.730 0.530 1.960 1.865 ;
        RECT  1.550 0.530 1.730 0.790 ;
        RECT  1.390 1.705 1.730 1.865 ;
        RECT  1.160 1.705 1.390 2.310 ;
        END
        AntennaDiffArea 0.406 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.275 0.505 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 -0.130 2.050 0.130 ;
        RECT  1.010 -0.130 1.270 0.695 ;
        RECT  0.330 -0.130 1.010 0.385 ;
        RECT  0.000 -0.130 0.330 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 2.740 2.050 3.000 ;
        RECT  1.655 2.050 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.100 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.980 1.365 1.550 1.525 ;
        RECT  0.820 0.890 0.980 1.920 ;
        RECT  0.700 0.890 0.820 1.050 ;
        RECT  0.370 1.760 0.820 1.920 ;
        RECT  0.540 0.635 0.700 1.050 ;
        RECT  0.440 0.635 0.540 0.895 ;
        RECT  0.140 1.760 0.370 2.100 ;
    END
END CLKBUFX3MTH

MACRO CLKBUFX40MTH
    CLASS CORE ;
    FOREIGN CLKBUFX40MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.145 0.425 9.315 1.610 ;
        RECT  8.995 0.425 9.145 2.395 ;
        RECT  8.885 0.900 8.995 2.395 ;
        RECT  8.235 0.900 8.885 1.980 ;
        RECT  7.915 0.425 8.235 2.485 ;
        RECT  7.295 0.900 7.915 1.980 ;
        RECT  6.975 0.425 7.295 2.485 ;
        RECT  6.325 0.900 6.975 1.980 ;
        RECT  6.215 0.900 6.325 2.485 ;
        RECT  6.065 0.415 6.215 2.485 ;
        RECT  5.895 0.415 6.065 1.980 ;
        RECT  5.245 0.900 5.895 1.980 ;
        RECT  4.040 0.430 5.245 2.485 ;
        RECT  2.965 0.430 4.040 0.910 ;
        RECT  3.105 1.545 4.040 2.485 ;
        END
        AntennaDiffArea 4.19 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.085 1.575 1.415 ;
        RECT  0.470 0.920 0.760 1.415 ;
        END
        AntennaGateArea 0.9347 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.745 -0.130 9.840 0.130 ;
        RECT  8.485 -0.130 8.745 0.680 ;
        RECT  6.725 -0.130 8.485 0.130 ;
        RECT  6.465 -0.130 6.725 0.680 ;
        RECT  4.705 -0.130 6.465 0.130 ;
        RECT  4.445 -0.130 4.705 0.250 ;
        RECT  2.685 -0.130 4.445 0.130 ;
        RECT  2.425 -0.130 2.685 0.695 ;
        RECT  1.605 -0.130 2.425 0.130 ;
        RECT  1.345 -0.130 1.605 0.300 ;
        RECT  0.525 -0.130 1.345 0.130 ;
        RECT  0.265 -0.130 0.525 0.695 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 2.740 9.840 3.000 ;
        RECT  9.425 1.805 9.685 3.000 ;
        RECT  5.785 2.740 9.425 3.000 ;
        RECT  5.525 2.230 5.785 3.000 ;
        RECT  0.925 2.740 5.525 3.000 ;
        RECT  0.665 2.225 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.405 1.095 3.735 1.295 ;
        RECT  2.145 1.095 2.405 2.315 ;
        RECT  1.885 0.435 2.145 1.295 ;
        RECT  1.465 1.715 2.145 2.005 ;
        RECT  1.065 0.485 1.885 0.695 ;
        RECT  1.205 1.715 1.465 2.315 ;
        RECT  0.385 1.715 1.205 2.005 ;
        RECT  0.805 0.435 1.065 0.695 ;
        RECT  0.125 1.715 0.385 2.315 ;
    END
END CLKBUFX40MTH

MACRO CLKBUFX4MTH
    CLASS CORE ;
    FOREIGN CLKBUFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.730 0.555 1.960 1.990 ;
        RECT  1.655 0.555 1.730 0.815 ;
        RECT  1.475 1.760 1.730 1.990 ;
        RECT  1.145 1.760 1.475 2.360 ;
        END
        AntennaDiffArea 0.541 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.595 1.580 ;
        END
        AntennaGateArea 0.0962 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.375 -0.130 2.050 0.130 ;
        RECT  1.115 -0.130 1.375 1.020 ;
        RECT  0.435 -0.130 1.115 0.515 ;
        RECT  0.000 -0.130 0.435 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 2.740 2.050 3.000 ;
        RECT  1.655 2.250 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.100 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.935 1.275 1.550 1.535 ;
        RECT  0.775 0.950 0.935 1.920 ;
        RECT  0.385 0.950 0.775 1.110 ;
        RECT  0.385 1.760 0.775 1.920 ;
        RECT  0.125 0.765 0.385 1.110 ;
        RECT  0.125 1.760 0.385 2.220 ;
    END
END CLKBUFX4MTH

MACRO CLKBUFX6MTH
    CLASS CORE ;
    FOREIGN CLKBUFX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 1.725 2.335 2.120 ;
        RECT  1.950 1.725 2.065 1.995 ;
        RECT  1.800 1.285 1.950 1.995 ;
        RECT  1.530 0.740 1.800 1.995 ;
        RECT  1.385 1.725 1.530 1.995 ;
        RECT  1.125 1.725 1.385 2.415 ;
        END
        AntennaDiffArea 0.718 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.255 0.555 1.580 ;
        END
        AntennaGateArea 0.1456 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  2.075 -0.130 2.335 1.025 ;
        RECT  1.635 -0.130 2.075 0.130 ;
        RECT  1.085 -0.130 1.635 0.300 ;
        RECT  0.825 -0.130 1.085 0.650 ;
        RECT  0.695 -0.130 0.825 0.300 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 2.740 2.460 3.000 ;
        RECT  1.665 2.570 2.265 3.000 ;
        RECT  0.000 2.740 1.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.945 1.205 1.215 1.465 ;
        RECT  0.785 0.865 0.945 1.920 ;
        RECT  0.385 0.865 0.785 1.025 ;
        RECT  0.385 1.760 0.785 1.920 ;
        RECT  0.125 0.765 0.385 1.025 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END CLKBUFX6MTH

MACRO CLKBUFX8MTH
    CLASS CORE ;
    FOREIGN CLKBUFX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.480 1.730 2.795 2.160 ;
        RECT  2.455 0.770 2.480 2.160 ;
        RECT  2.050 0.770 2.455 2.070 ;
        RECT  1.775 0.770 2.050 1.110 ;
        RECT  1.770 1.730 2.050 2.070 ;
        RECT  1.435 0.595 1.775 1.110 ;
        RECT  1.430 1.730 1.770 2.400 ;
        END
        AntennaDiffArea 0.861 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.245 0.855 1.505 ;
        RECT  0.100 1.245 0.310 1.580 ;
        END
        AntennaGateArea 0.1963 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.130 3.280 0.130 ;
        RECT  2.525 -0.130 3.125 0.590 ;
        RECT  2.275 -0.130 2.525 0.130 ;
        RECT  2.015 -0.130 2.275 0.590 ;
        RECT  1.190 -0.130 2.015 0.130 ;
        RECT  0.930 -0.130 1.190 0.710 ;
        RECT  0.740 -0.130 0.930 0.130 ;
        RECT  0.140 -0.130 0.740 0.380 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.895 2.570 3.155 3.000 ;
        RECT  2.245 2.740 2.895 3.000 ;
        RECT  1.985 2.255 2.245 3.000 ;
        RECT  1.175 2.740 1.985 3.000 ;
        RECT  0.235 2.495 1.175 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.225 1.290 1.665 1.550 ;
        RECT  1.065 0.905 1.225 1.850 ;
        RECT  0.650 0.905 1.065 1.065 ;
        RECT  0.790 1.690 1.065 1.850 ;
        RECT  0.530 1.690 0.790 2.070 ;
        RECT  0.390 0.740 0.650 1.065 ;
    END
END CLKBUFX8MTH

MACRO CLKINVX12MTH
    CLASS CORE ;
    FOREIGN CLKINVX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.650 1.800 2.755 2.400 ;
        RECT  2.495 0.680 2.650 2.400 ;
        RECT  2.390 0.680 2.495 2.200 ;
        RECT  1.940 0.770 2.390 2.200 ;
        RECT  1.540 0.770 1.940 1.090 ;
        RECT  1.825 1.800 1.940 2.200 ;
        RECT  1.565 1.800 1.825 2.400 ;
        RECT  0.895 1.800 1.565 2.200 ;
        RECT  1.220 0.390 1.540 1.090 ;
        RECT  0.635 1.800 0.895 2.400 ;
        END
        AntennaDiffArea 1.431 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.290 1.745 1.580 ;
        END
        AntennaGateArea 0.9295 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.105 -0.130 3.280 0.130 ;
        RECT  2.265 -0.130 3.105 0.435 ;
        RECT  2.080 -0.130 2.265 0.130 ;
        RECT  1.820 -0.130 2.080 0.590 ;
        RECT  0.940 -0.130 1.820 0.130 ;
        RECT  0.340 -0.130 0.940 0.995 ;
        RECT  0.000 -0.130 0.340 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 3.280 3.000 ;
        RECT  0.125 1.875 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX12MTH

MACRO CLKINVX16MTH
    CLASS CORE ;
    FOREIGN CLKINVX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.715 1.565 3.975 2.400 ;
        RECT  3.240 1.565 3.715 2.095 ;
        RECT  2.955 0.435 3.240 2.095 ;
        RECT  2.695 0.435 2.955 2.400 ;
        RECT  2.355 0.435 2.695 2.095 ;
        RECT  0.670 0.435 2.355 0.955 ;
        RECT  1.935 1.565 2.355 2.095 ;
        RECT  1.675 1.565 1.935 2.400 ;
        RECT  0.930 1.565 1.675 2.095 ;
        RECT  0.670 1.565 0.930 2.400 ;
        END
        AntennaDiffArea 2.019 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.175 2.120 1.335 ;
        RECT  0.100 1.175 0.310 1.580 ;
        END
        AntennaGateArea 1.2363 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.810 -0.130 4.100 0.130 ;
        RECT  3.550 -0.130 3.810 0.640 ;
        RECT  2.670 -0.130 3.550 0.130 ;
        RECT  2.410 -0.130 2.670 0.250 ;
        RECT  1.530 -0.130 2.410 0.130 ;
        RECT  1.270 -0.130 1.530 0.250 ;
        RECT  0.390 -0.130 1.270 0.130 ;
        RECT  0.130 -0.130 0.390 0.640 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 2.740 4.100 3.000 ;
        RECT  3.205 2.305 3.465 3.000 ;
        RECT  2.445 2.740 3.205 3.000 ;
        RECT  2.185 2.305 2.445 3.000 ;
        RECT  0.385 2.740 2.185 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX16MTH

MACRO CLKINVX1MTH
    CLASS CORE ;
    FOREIGN CLKINVX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.760 1.130 2.020 ;
        RECT  0.710 0.760 0.920 1.020 ;
        RECT  0.680 1.760 0.920 2.020 ;
        END
        AntennaDiffArea 0.276 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.225 1.240 0.720 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 -0.130 1.230 0.130 ;
        RECT  0.690 -0.130 0.950 0.510 ;
        RECT  0.400 -0.130 0.690 0.130 ;
        RECT  0.140 -0.130 0.400 1.020 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.940 2.740 1.230 3.000 ;
        RECT  0.680 2.495 0.940 3.000 ;
        RECT  0.400 2.740 0.680 3.000 ;
        RECT  0.140 1.825 0.400 3.000 ;
        RECT  0.000 2.740 0.140 3.000 ;
        END
    END VDD
END CLKINVX1MTH

MACRO CLKINVX20MTH
    CLASS CORE ;
    FOREIGN CLKINVX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 0.435 3.875 2.420 ;
        RECT  2.865 0.435 3.565 2.325 ;
        RECT  2.605 0.435 2.865 2.425 ;
        RECT  0.665 0.435 2.605 0.835 ;
        RECT  1.895 1.485 2.605 2.325 ;
        RECT  1.635 1.485 1.895 2.425 ;
        RECT  0.925 1.485 1.635 2.325 ;
        RECT  0.665 1.485 0.925 2.400 ;
        END
        AntennaDiffArea 2.338 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.055 2.290 1.215 ;
        RECT  0.100 1.055 0.310 1.580 ;
        END
        AntennaGateArea 1.5457 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  4.125 -0.130 4.385 0.670 ;
        RECT  2.405 -0.130 4.125 0.130 ;
        RECT  2.145 -0.130 2.405 0.250 ;
        RECT  0.385 -0.130 2.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.675 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.890 4.385 3.000 ;
        RECT  0.385 2.740 4.125 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX20MTH

MACRO CLKINVX24MTH
    CLASS CORE ;
    FOREIGN CLKINVX24MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.440 1.160 4.700 2.440 ;
        RECT  3.835 1.760 4.440 2.160 ;
        RECT  3.745 0.755 3.835 2.160 ;
        RECT  3.485 0.755 3.745 2.400 ;
        RECT  3.135 0.755 3.485 2.160 ;
        RECT  2.940 0.755 3.135 1.085 ;
        RECT  2.805 1.760 3.135 2.160 ;
        RECT  2.680 0.465 2.940 1.085 ;
        RECT  2.545 1.760 2.805 2.400 ;
        RECT  1.920 0.755 2.680 1.085 ;
        RECT  1.855 1.760 2.545 2.160 ;
        RECT  1.660 0.425 1.920 1.085 ;
        RECT  1.595 1.760 1.855 2.400 ;
        RECT  0.900 0.755 1.660 1.085 ;
        RECT  0.925 1.760 1.595 2.160 ;
        RECT  0.665 1.760 0.925 2.400 ;
        RECT  0.640 0.425 0.900 1.085 ;
        END
        AntennaDiffArea 2.7 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.305 2.770 1.540 ;
        END
        AntennaGateArea 1.8486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.565 -0.130 5.740 0.130 ;
        RECT  4.965 -0.130 5.565 0.300 ;
        RECT  4.695 -0.130 4.965 0.130 ;
        RECT  3.755 -0.130 4.695 0.300 ;
        RECT  3.480 -0.130 3.755 0.130 ;
        RECT  3.220 -0.130 3.480 0.300 ;
        RECT  2.430 -0.130 3.220 0.130 ;
        RECT  2.170 -0.130 2.430 0.565 ;
        RECT  1.410 -0.130 2.170 0.130 ;
        RECT  1.150 -0.130 1.410 0.565 ;
        RECT  0.390 -0.130 1.150 0.130 ;
        RECT  0.130 -0.130 0.390 0.990 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.580 2.740 5.740 3.000 ;
        RECT  4.980 1.685 5.580 3.000 ;
        RECT  0.385 2.740 4.980 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX24MTH

MACRO CLKINVX2MTH
    CLASS CORE ;
    FOREIGN CLKINVX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.755 1.130 2.360 ;
        RECT  0.740 0.755 0.920 1.015 ;
        RECT  0.740 1.760 0.920 2.360 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.195 0.720 1.580 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.970 -0.130 1.230 0.130 ;
        RECT  0.710 -0.130 0.970 0.445 ;
        RECT  0.460 -0.130 0.710 0.130 ;
        RECT  0.200 -0.130 0.460 1.005 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 2.740 1.230 3.000 ;
        RECT  0.200 1.850 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
END CLKINVX2MTH

MACRO CLKINVX32MTH
    CLASS CORE ;
    FOREIGN CLKINVX32MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.520 0.745 6.840 2.365 ;
        RECT  5.825 0.745 6.520 1.535 ;
        RECT  5.565 0.745 5.825 2.475 ;
        RECT  4.820 0.745 5.565 1.535 ;
        RECT  4.540 0.745 4.820 2.410 ;
        RECT  3.870 0.745 4.540 1.535 ;
        RECT  3.590 0.745 3.870 2.370 ;
        RECT  3.445 0.745 3.590 1.535 ;
        RECT  3.185 0.425 3.445 1.535 ;
        RECT  3.075 0.745 3.185 1.535 ;
        RECT  2.675 0.745 3.075 2.365 ;
        RECT  2.425 0.745 2.675 2.120 ;
        RECT  2.165 0.385 2.425 2.120 ;
        RECT  1.995 0.745 2.165 2.120 ;
        RECT  1.405 0.745 1.995 1.075 ;
        RECT  1.915 1.760 1.995 2.120 ;
        RECT  1.655 1.760 1.915 2.365 ;
        RECT  0.895 1.760 1.655 2.120 ;
        RECT  1.145 0.385 1.405 1.075 ;
        RECT  0.385 0.745 1.145 1.075 ;
        RECT  0.635 1.760 0.895 2.365 ;
        RECT  0.125 0.395 0.385 1.075 ;
        END
        AntennaDiffArea 3.875 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.295 1.745 1.540 ;
        END
        AntennaGateArea 2.4479 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 -0.130 6.970 0.130 ;
        RECT  3.725 -0.130 3.985 0.565 ;
        RECT  2.935 -0.130 3.725 0.130 ;
        RECT  2.675 -0.130 2.935 0.565 ;
        RECT  1.915 -0.130 2.675 0.130 ;
        RECT  1.655 -0.130 1.915 0.565 ;
        RECT  0.895 -0.130 1.655 0.130 ;
        RECT  0.635 -0.130 0.895 0.565 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 2.740 6.970 3.000 ;
        RECT  6.075 1.830 6.335 3.000 ;
        RECT  5.315 2.740 6.075 3.000 ;
        RECT  5.055 1.850 5.315 3.000 ;
        RECT  2.425 2.740 5.055 3.000 ;
        RECT  2.165 2.305 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 2.305 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.870 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX32MTH

MACRO CLKINVX3MTH
    CLASS CORE ;
    FOREIGN CLKINVX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 0.710 1.150 1.990 ;
        RECT  0.920 0.710 0.925 2.260 ;
        RECT  0.665 0.710 0.920 0.970 ;
        RECT  0.665 1.760 0.920 2.260 ;
        END
        AntennaDiffArea 0.406 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 1.160 0.720 1.580 ;
        END
        AntennaGateArea 0.2314 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 -0.130 1.640 0.130 ;
        RECT  0.730 -0.130 1.330 0.315 ;
        RECT  0.385 -0.130 0.730 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 2.740 1.640 3.000 ;
        RECT  1.205 2.170 1.465 3.000 ;
        RECT  0.385 2.740 1.205 3.000 ;
        RECT  0.125 1.780 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX3MTH

MACRO CLKINVX40MTH
    CLASS CORE ;
    FOREIGN CLKINVX40MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.685 0.875 7.945 2.420 ;
        RECT  7.405 0.875 7.685 1.955 ;
        RECT  7.145 0.430 7.405 1.955 ;
        RECT  6.965 0.875 7.145 1.955 ;
        RECT  6.705 0.875 6.965 2.470 ;
        RECT  6.325 0.875 6.705 1.955 ;
        RECT  6.065 0.430 6.325 1.955 ;
        RECT  5.945 0.875 6.065 1.955 ;
        RECT  5.685 0.875 5.945 2.470 ;
        RECT  5.245 0.875 5.685 1.955 ;
        RECT  4.985 0.430 5.245 1.955 ;
        RECT  4.975 0.875 4.985 1.955 ;
        RECT  4.715 0.875 4.975 2.470 ;
        RECT  4.165 0.875 4.715 1.955 ;
        RECT  3.905 0.430 4.165 1.955 ;
        RECT  3.895 0.875 3.905 1.955 ;
        RECT  3.635 0.875 3.895 2.470 ;
        RECT  3.085 0.875 3.635 1.955 ;
        RECT  2.925 0.430 3.085 1.955 ;
        RECT  2.665 0.430 2.925 2.420 ;
        RECT  1.905 0.430 2.665 2.120 ;
        RECT  1.785 0.430 1.905 2.420 ;
        RECT  0.665 0.430 1.785 0.900 ;
        RECT  1.205 1.420 1.785 2.420 ;
        RECT  0.665 1.720 1.205 2.420 ;
        END
        AntennaDiffArea 4.543 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.080 1.605 1.240 ;
        RECT  0.470 1.080 0.760 1.540 ;
        END
        AntennaGateArea 3.0628 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.315 -0.130 8.610 0.130 ;
        RECT  7.715 -0.130 8.315 0.695 ;
        RECT  6.865 -0.130 7.715 0.130 ;
        RECT  6.605 -0.130 6.865 0.695 ;
        RECT  5.785 -0.130 6.605 0.130 ;
        RECT  5.525 -0.130 5.785 0.695 ;
        RECT  4.705 -0.130 5.525 0.130 ;
        RECT  4.445 -0.130 4.705 0.695 ;
        RECT  3.625 -0.130 4.445 0.130 ;
        RECT  3.365 -0.130 3.625 0.695 ;
        RECT  2.545 -0.130 3.365 0.130 ;
        RECT  2.285 -0.130 2.545 0.250 ;
        RECT  1.465 -0.130 2.285 0.130 ;
        RECT  1.205 -0.130 1.465 0.250 ;
        RECT  0.385 -0.130 1.205 0.130 ;
        RECT  0.125 -0.130 0.385 0.715 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.485 2.740 8.610 3.000 ;
        RECT  8.225 1.755 8.485 3.000 ;
        RECT  6.455 2.740 8.225 3.000 ;
        RECT  6.195 2.140 6.455 3.000 ;
        RECT  4.435 2.740 6.195 3.000 ;
        RECT  4.175 2.225 4.435 3.000 ;
        RECT  2.415 2.740 4.175 3.000 ;
        RECT  2.155 2.300 2.415 3.000 ;
        RECT  0.385 2.740 2.155 3.000 ;
        RECT  0.125 1.820 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX40MTH

MACRO CLKINVX4MTH
    CLASS CORE ;
    FOREIGN CLKINVX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 0.425 1.390 1.025 ;
        RECT  1.040 0.425 1.270 2.010 ;
        RECT  0.950 1.700 1.040 2.010 ;
        RECT  0.920 1.700 0.950 2.380 ;
        RECT  0.690 1.780 0.920 2.380 ;
        END
        AntennaDiffArea 0.583 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.275 0.730 1.580 ;
        END
        AntennaGateArea 0.3068 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.820 -0.130 1.640 0.130 ;
        RECT  0.220 -0.130 0.820 1.025 ;
        RECT  0.000 -0.130 0.220 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.490 2.740 1.640 3.000 ;
        RECT  1.230 2.245 1.490 3.000 ;
        RECT  0.410 2.740 1.230 3.000 ;
        RECT  0.150 1.890 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
END CLKINVX4MTH

MACRO CLKINVX6MTH
    CLASS CORE ;
    FOREIGN CLKINVX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 1.730 1.915 2.380 ;
        RECT  1.505 1.730 1.655 1.990 ;
        RECT  1.245 0.850 1.505 1.990 ;
        RECT  1.190 0.850 1.245 1.110 ;
        RECT  0.895 1.730 1.245 1.990 ;
        RECT  0.930 0.680 1.190 1.110 ;
        RECT  0.635 1.730 0.895 2.380 ;
        END
        AntennaDiffArea 0.8 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.290 1.065 1.550 ;
        END
        AntennaGateArea 0.4589 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.730 -0.130 2.050 0.130 ;
        RECT  1.470 -0.130 1.730 0.670 ;
        RECT  0.650 -0.130 1.470 0.130 ;
        RECT  0.390 -0.130 0.650 1.025 ;
        RECT  0.000 -0.130 0.390 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 2.740 2.050 3.000 ;
        RECT  1.145 2.200 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.915 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX6MTH

MACRO CLKINVX8MTH
    CLASS CORE ;
    FOREIGN CLKINVX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 1.730 1.825 2.330 ;
        RECT  1.295 0.425 1.635 2.330 ;
        RECT  0.895 1.730 1.295 2.030 ;
        RECT  0.635 1.730 0.895 2.330 ;
        END
        AntennaDiffArea 0.956 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.290 1.065 1.550 ;
        END
        AntennaGateArea 0.6136 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.125 -0.130 2.460 0.130 ;
        RECT  1.865 -0.130 2.125 1.025 ;
        RECT  0.905 -0.130 1.865 0.130 ;
        RECT  0.305 -0.130 0.905 1.025 ;
        RECT  0.000 -0.130 0.305 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  2.075 1.840 2.335 3.000 ;
        RECT  0.385 2.740 2.075 3.000 ;
        RECT  0.125 1.855 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKINVX8MTH

MACRO CLKMX2X12MTH
    CLASS CORE ;
    FOREIGN CLKMX2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 0.715 6.020 2.435 ;
        RECT  5.140 0.715 5.760 1.335 ;
        RECT  5.000 0.455 5.140 1.335 ;
        RECT  4.800 0.455 5.000 2.455 ;
        RECT  4.740 0.715 4.800 2.455 ;
        RECT  3.980 0.715 4.740 1.335 ;
        RECT  3.720 0.440 3.980 2.455 ;
        END
        AntennaDiffArea 1.48 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.430 1.205 0.720 1.700 ;
        END
        AntennaGateArea 0.2288 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.070 1.520 1.130 1.990 ;
        RECT  0.910 1.230 1.070 1.990 ;
        END
        AntennaGateArea 0.1534 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.830 1.120 3.180 1.580 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.940 -0.130 6.150 0.130 ;
        RECT  5.340 -0.130 5.940 0.535 ;
        RECT  4.520 -0.130 5.340 0.130 ;
        RECT  4.260 -0.130 4.520 0.535 ;
        RECT  3.440 -0.130 4.260 0.130 ;
        RECT  3.180 -0.130 3.440 0.690 ;
        RECT  0.955 -0.130 3.180 0.130 ;
        RECT  0.690 -0.130 0.955 0.685 ;
        RECT  0.385 -0.130 0.690 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.510 2.740 6.150 3.000 ;
        RECT  5.250 1.835 5.510 3.000 ;
        RECT  4.490 2.740 5.250 3.000 ;
        RECT  4.230 1.575 4.490 3.000 ;
        RECT  3.430 2.740 4.230 3.000 ;
        RECT  3.170 2.100 3.430 3.000 ;
        RECT  0.925 2.740 3.170 3.000 ;
        RECT  0.665 2.175 0.925 3.000 ;
        RECT  0.295 2.570 0.665 3.000 ;
        RECT  0.000 2.740 0.295 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.365 0.980 3.525 1.920 ;
        RECT  2.990 1.760 3.365 1.920 ;
        RECT  2.830 1.760 2.990 2.385 ;
        RECT  2.665 0.510 2.875 0.825 ;
        RECT  2.265 2.225 2.830 2.385 ;
        RECT  2.650 0.665 2.665 0.825 ;
        RECT  2.490 0.665 2.650 2.005 ;
        RECT  1.410 0.310 2.485 0.470 ;
        RECT  2.105 0.665 2.265 2.385 ;
        RECT  1.685 2.125 2.105 2.385 ;
        RECT  1.765 0.655 1.925 1.765 ;
        RECT  1.590 0.655 1.765 0.915 ;
        RECT  1.495 1.605 1.765 1.765 ;
        RECT  1.410 1.125 1.585 1.385 ;
        RECT  1.335 1.605 1.495 2.405 ;
        RECT  1.250 0.310 1.410 1.385 ;
        RECT  1.175 2.175 1.335 2.405 ;
        RECT  0.385 0.865 1.250 1.025 ;
        RECT  0.250 0.665 0.385 1.025 ;
        RECT  0.250 1.895 0.385 2.155 ;
        RECT  0.090 0.665 0.250 2.155 ;
    END
END CLKMX2X12MTH

MACRO CLKMX2X16MTH
    CLASS CORE ;
    FOREIGN CLKMX2X16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.465 0.385 6.835 1.785 ;
        RECT  6.305 1.085 6.465 1.785 ;
        RECT  6.045 1.085 6.305 2.325 ;
        RECT  5.825 1.085 6.045 1.785 ;
        RECT  5.325 0.430 5.825 1.785 ;
        RECT  4.945 0.430 5.325 2.440 ;
        RECT  3.555 0.430 4.945 0.810 ;
        RECT  3.885 2.060 4.945 2.440 ;
        END
        AntennaDiffArea 1.862 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 2.275 1.835 2.540 ;
        RECT  0.770 2.275 1.575 2.435 ;
        RECT  0.555 2.110 0.770 2.435 ;
        RECT  0.295 2.110 0.555 2.475 ;
        RECT  0.245 2.315 0.295 2.475 ;
        END
        AntennaGateArea 0.2288 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.675 0.905 1.205 1.170 ;
        END
        AntennaGateArea 0.1534 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 1.330 3.630 1.540 ;
        RECT  2.955 1.330 3.180 1.490 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.285 -0.130 6.970 0.130 ;
        RECT  6.075 -0.130 6.285 0.670 ;
        RECT  4.355 -0.130 6.075 0.130 ;
        RECT  4.095 -0.130 4.355 0.250 ;
        RECT  1.005 -0.130 4.095 0.130 ;
        RECT  0.745 -0.130 1.005 0.660 ;
        RECT  0.345 -0.130 0.745 0.320 ;
        RECT  0.000 -0.130 0.345 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 2.065 6.845 3.000 ;
        RECT  5.765 2.740 6.585 3.000 ;
        RECT  5.505 2.065 5.765 3.000 ;
        RECT  4.685 2.740 5.505 3.000 ;
        RECT  4.425 2.620 4.685 3.000 ;
        RECT  3.600 2.740 4.425 3.000 ;
        RECT  3.340 2.510 3.600 3.000 ;
        RECT  0.925 2.740 3.340 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.970 0.990 4.545 1.245 ;
        RECT  3.810 0.990 3.970 1.880 ;
        RECT  3.115 0.990 3.810 1.150 ;
        RECT  3.460 1.720 3.810 1.880 ;
        RECT  3.300 1.720 3.460 2.330 ;
        RECT  2.545 2.170 3.300 2.330 ;
        RECT  2.955 0.310 3.115 1.150 ;
        RECT  2.795 1.670 3.055 1.970 ;
        RECT  2.055 0.310 2.955 0.470 ;
        RECT  2.775 1.670 2.795 1.830 ;
        RECT  2.615 0.650 2.775 1.830 ;
        RECT  2.285 2.005 2.545 2.330 ;
        RECT  2.275 0.840 2.435 1.785 ;
        RECT  1.545 0.840 2.275 1.000 ;
        RECT  2.060 1.625 2.275 1.785 ;
        RECT  1.935 1.185 2.095 1.445 ;
        RECT  1.900 1.625 2.060 1.905 ;
        RECT  1.795 0.310 2.055 0.615 ;
        RECT  1.565 1.285 1.935 1.445 ;
        RECT  1.465 1.745 1.900 1.905 ;
        RECT  1.405 1.285 1.565 1.510 ;
        RECT  1.385 0.415 1.545 1.000 ;
        RECT  1.205 1.745 1.465 2.020 ;
        RECT  0.385 1.350 1.405 1.510 ;
        RECT  1.285 0.415 1.385 0.675 ;
        RECT  0.335 0.590 0.435 0.850 ;
        RECT  0.335 1.350 0.385 1.920 ;
        RECT  0.175 0.590 0.335 1.920 ;
        RECT  0.125 1.760 0.175 1.920 ;
    END
END CLKMX2X16MTH

MACRO CLKMX2X2MTH
    CLASS CORE ;
    FOREIGN CLKMX2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.635 4.000 2.425 ;
        RECT  3.725 0.635 3.790 0.895 ;
        RECT  3.715 2.165 3.790 2.425 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.130 0.380 1.580 ;
        END
        AntennaGateArea 0.2132 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.185 1.375 ;
        END
        AntennaGateArea 0.1235 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.810 1.290 3.205 1.680 ;
        END
        AntennaGateArea 0.1235 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.905 -0.130 4.100 0.130 ;
        RECT  3.645 -0.130 3.905 0.300 ;
        RECT  3.405 -0.130 3.645 0.130 ;
        RECT  3.185 -0.130 3.405 0.770 ;
        RECT  0.955 -0.130 3.185 0.130 ;
        RECT  0.695 -0.130 0.955 0.575 ;
        RECT  0.385 -0.130 0.695 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.390 2.740 4.100 3.000 ;
        RECT  3.130 2.230 3.390 3.000 ;
        RECT  1.000 2.740 3.130 3.000 ;
        RECT  0.740 2.185 1.000 3.000 ;
        RECT  0.385 2.740 0.740 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.385 0.950 3.545 2.020 ;
        RECT  3.005 0.950 3.385 1.110 ;
        RECT  2.950 1.860 3.385 2.020 ;
        RECT  2.845 0.310 3.005 1.110 ;
        RECT  2.790 1.860 2.950 2.435 ;
        RECT  2.095 0.310 2.845 0.470 ;
        RECT  1.890 2.275 2.790 2.435 ;
        RECT  2.525 0.685 2.665 0.845 ;
        RECT  2.525 1.835 2.610 2.095 ;
        RECT  2.365 0.685 2.525 2.095 ;
        RECT  1.945 0.845 2.105 2.095 ;
        RECT  1.835 0.310 2.095 0.665 ;
        RECT  1.525 0.845 1.945 1.005 ;
        RECT  1.320 1.935 1.945 2.095 ;
        RECT  1.605 1.185 1.765 1.755 ;
        RECT  0.740 1.595 1.605 1.755 ;
        RECT  1.365 0.540 1.525 1.005 ;
        RECT  1.265 0.540 1.365 0.700 ;
        RECT  0.560 0.755 0.740 2.005 ;
        RECT  0.385 0.755 0.560 0.915 ;
        RECT  0.385 1.845 0.560 2.005 ;
        RECT  0.125 0.685 0.385 0.915 ;
        RECT  0.125 1.845 0.385 2.105 ;
    END
END CLKMX2X2MTH

MACRO CLKMX2X3MTH
    CLASS CORE ;
    FOREIGN CLKMX2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.225 1.290 4.410 1.580 ;
        RECT  4.065 0.745 4.225 1.795 ;
        RECT  3.965 0.745 4.065 1.005 ;
        RECT  3.945 1.635 4.065 1.795 ;
        RECT  3.785 1.635 3.945 2.230 ;
        RECT  3.615 2.070 3.785 2.230 ;
        END
        AntennaDiffArea 0.458 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.480 2.230 1.740 2.560 ;
        RECT  0.760 2.230 1.480 2.390 ;
        RECT  0.245 2.150 0.760 2.475 ;
        END
        AntennaGateArea 0.2288 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 0.890 1.170 1.365 ;
        END
        AntennaGateArea 0.1547 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.110 3.220 1.540 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.225 -0.130 4.510 0.130 ;
        RECT  3.425 -0.130 4.225 0.300 ;
        RECT  0.955 -0.130 3.425 0.130 ;
        RECT  0.355 -0.130 0.955 0.300 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.995 4.385 3.000 ;
        RECT  1.300 2.740 4.125 3.000 ;
        RECT  1.080 2.570 1.300 3.000 ;
        RECT  0.000 2.740 1.080 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.560 1.185 3.880 1.455 ;
        RECT  3.410 0.535 3.560 1.880 ;
        RECT  3.400 0.535 3.410 2.355 ;
        RECT  3.220 0.535 3.400 0.695 ;
        RECT  3.250 1.720 3.400 2.355 ;
        RECT  2.175 2.195 3.250 2.355 ;
        RECT  3.060 0.315 3.220 0.695 ;
        RECT  2.065 0.315 3.060 0.475 ;
        RECT  2.750 1.850 2.945 2.010 ;
        RECT  2.750 0.655 2.875 0.815 ;
        RECT  2.590 0.655 2.750 2.010 ;
        RECT  2.250 0.770 2.410 1.975 ;
        RECT  1.510 0.770 2.250 0.930 ;
        RECT  1.895 1.815 2.250 1.975 ;
        RECT  1.910 1.125 2.070 1.560 ;
        RECT  1.795 0.315 2.065 0.590 ;
        RECT  1.535 1.400 1.910 1.560 ;
        RECT  1.720 1.815 1.895 2.045 ;
        RECT  1.065 1.885 1.720 2.045 ;
        RECT  1.375 1.400 1.535 1.705 ;
        RECT  1.350 0.550 1.510 0.930 ;
        RECT  0.385 1.545 1.375 1.705 ;
        RECT  1.235 0.550 1.350 0.710 ;
        RECT  0.225 0.560 0.385 1.970 ;
        RECT  0.125 0.560 0.225 0.820 ;
        RECT  0.125 1.710 0.225 1.970 ;
    END
END CLKMX2X3MTH

MACRO CLKMX2X4MTH
    CLASS CORE ;
    FOREIGN CLKMX2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.150 0.575 4.410 1.785 ;
        RECT  3.995 0.575 4.150 0.835 ;
        RECT  3.945 1.625 4.150 1.785 ;
        RECT  3.785 1.625 3.945 2.365 ;
        RECT  3.615 2.105 3.785 2.365 ;
        END
        AntennaDiffArea 0.559 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.480 2.230 1.740 2.560 ;
        RECT  0.720 2.230 1.480 2.390 ;
        RECT  0.245 2.110 0.720 2.475 ;
        END
        AntennaGateArea 0.2288 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 0.880 1.155 1.360 ;
        END
        AntennaGateArea 0.1547 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 0.995 3.180 1.580 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.685 -0.130 4.510 0.130 ;
        RECT  3.425 -0.130 3.685 0.300 ;
        RECT  0.955 -0.130 3.425 0.130 ;
        RECT  0.355 -0.130 0.955 0.300 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.965 4.385 3.000 ;
        RECT  1.300 2.740 4.125 3.000 ;
        RECT  1.080 2.570 1.300 3.000 ;
        RECT  0.000 2.740 1.080 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.605 1.185 3.880 1.445 ;
        RECT  3.445 0.550 3.605 1.920 ;
        RECT  3.245 0.550 3.445 0.710 ;
        RECT  3.285 1.760 3.445 1.920 ;
        RECT  3.125 1.760 3.285 2.355 ;
        RECT  3.085 0.315 3.245 0.710 ;
        RECT  2.175 2.195 3.125 2.355 ;
        RECT  2.055 0.315 3.085 0.475 ;
        RECT  2.775 1.760 2.945 1.920 ;
        RECT  2.775 0.655 2.875 0.815 ;
        RECT  2.615 0.655 2.775 1.920 ;
        RECT  2.275 0.770 2.435 1.970 ;
        RECT  1.615 0.770 2.275 0.930 ;
        RECT  1.895 1.810 2.275 1.970 ;
        RECT  1.935 1.125 2.095 1.620 ;
        RECT  1.795 0.315 2.055 0.590 ;
        RECT  1.495 1.460 1.935 1.620 ;
        RECT  1.730 1.810 1.895 2.045 ;
        RECT  1.065 1.885 1.730 2.045 ;
        RECT  1.455 0.540 1.615 0.930 ;
        RECT  1.335 1.460 1.495 1.705 ;
        RECT  1.170 0.540 1.455 0.700 ;
        RECT  0.385 1.545 1.335 1.705 ;
        RECT  0.225 0.610 0.385 1.920 ;
        RECT  0.125 0.610 0.225 0.770 ;
        RECT  0.125 1.760 0.225 1.920 ;
    END
END CLKMX2X4MTH

MACRO CLKMX2X6MTH
    CLASS CORE ;
    FOREIGN CLKMX2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 1.625 5.205 2.360 ;
        RECT  4.860 1.625 4.945 1.785 ;
        RECT  4.570 0.835 4.860 1.785 ;
        RECT  4.320 0.835 4.570 0.995 ;
        RECT  4.255 1.625 4.570 1.785 ;
        RECT  4.060 0.575 4.320 0.995 ;
        RECT  4.095 1.625 4.255 2.465 ;
        RECT  3.905 2.205 4.095 2.465 ;
        END
        AntennaDiffArea 0.839 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 2.275 1.835 2.540 ;
        RECT  0.760 2.275 1.575 2.435 ;
        RECT  0.505 2.150 0.760 2.435 ;
        RECT  0.245 2.150 0.505 2.475 ;
        END
        AntennaGateArea 0.2288 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.295 1.405 ;
        END
        AntennaGateArea 0.1547 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.030 3.295 1.580 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.200 -0.130 5.330 0.130 ;
        RECT  4.600 -0.130 5.200 0.655 ;
        RECT  3.680 -0.130 4.600 0.130 ;
        RECT  3.420 -0.130 3.680 0.360 ;
        RECT  0.965 -0.130 3.420 0.130 ;
        RECT  0.705 -0.130 0.965 0.700 ;
        RECT  0.000 -0.130 0.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.695 2.740 5.330 3.000 ;
        RECT  4.435 1.965 4.695 3.000 ;
        RECT  3.625 2.740 4.435 3.000 ;
        RECT  3.365 2.570 3.625 3.000 ;
        RECT  0.925 2.740 3.365 3.000 ;
        RECT  0.665 2.615 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.855 1.180 4.335 1.440 ;
        RECT  3.695 0.540 3.855 2.025 ;
        RECT  3.240 0.540 3.695 0.700 ;
        RECT  3.445 1.865 3.695 2.025 ;
        RECT  3.285 1.865 3.445 2.355 ;
        RECT  2.315 2.195 3.285 2.355 ;
        RECT  3.080 0.315 3.240 0.700 ;
        RECT  2.790 1.760 3.085 1.920 ;
        RECT  2.095 0.315 3.080 0.475 ;
        RECT  2.790 0.655 2.895 0.815 ;
        RECT  2.630 0.655 2.790 1.920 ;
        RECT  2.290 0.770 2.450 1.975 ;
        RECT  1.635 0.770 2.290 0.930 ;
        RECT  2.035 1.815 2.290 1.975 ;
        RECT  1.950 1.125 2.110 1.635 ;
        RECT  1.835 0.315 2.095 0.590 ;
        RECT  1.850 1.815 2.035 2.090 ;
        RECT  1.625 1.475 1.950 1.635 ;
        RECT  1.205 1.930 1.850 2.090 ;
        RECT  1.475 0.540 1.635 0.930 ;
        RECT  1.465 1.475 1.625 1.750 ;
        RECT  1.255 0.540 1.475 0.700 ;
        RECT  0.385 1.590 1.465 1.750 ;
        RECT  0.225 0.500 0.385 1.970 ;
        RECT  0.125 0.500 0.225 0.760 ;
        RECT  0.125 1.710 0.225 1.970 ;
    END
END CLKMX2X6MTH

MACRO CLKMX2X8MTH
    CLASS CORE ;
    FOREIGN CLKMX2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 0.845 5.235 1.795 ;
        RECT  4.815 0.845 5.075 2.360 ;
        RECT  4.285 0.845 4.815 1.005 ;
        RECT  4.335 1.635 4.815 1.795 ;
        RECT  4.175 1.635 4.335 1.950 ;
        RECT  4.125 0.575 4.285 1.005 ;
        RECT  4.075 1.790 4.175 1.950 ;
        RECT  4.010 0.575 4.125 0.835 ;
        RECT  3.815 1.790 4.075 2.390 ;
        END
        AntennaDiffArea 0.896 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 2.275 1.835 2.540 ;
        RECT  0.720 2.275 1.575 2.435 ;
        RECT  0.505 2.110 0.720 2.435 ;
        RECT  0.245 2.110 0.505 2.475 ;
        END
        AntennaGateArea 0.2288 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 0.880 1.225 1.405 ;
        END
        AntennaGateArea 0.1534 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.110 3.270 1.580 ;
        END
        AntennaGateArea 0.1534 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 -0.130 5.740 0.130 ;
        RECT  4.550 -0.130 5.150 0.660 ;
        RECT  3.730 -0.130 4.550 0.130 ;
        RECT  3.470 -0.130 3.730 0.590 ;
        RECT  0.955 -0.130 3.470 0.130 ;
        RECT  0.695 -0.130 0.955 0.700 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 1.965 5.615 3.000 ;
        RECT  0.925 2.740 5.355 3.000 ;
        RECT  0.665 2.620 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.610 1.185 4.590 1.455 ;
        RECT  3.450 0.770 3.610 2.355 ;
        RECT  3.290 0.770 3.450 0.930 ;
        RECT  2.315 2.195 3.450 2.355 ;
        RECT  3.130 0.315 3.290 0.930 ;
        RECT  2.055 0.315 3.130 0.475 ;
        RECT  2.775 1.760 3.085 1.920 ;
        RECT  2.775 0.655 2.945 0.815 ;
        RECT  2.615 0.655 2.775 1.920 ;
        RECT  2.275 0.770 2.435 1.975 ;
        RECT  1.615 0.770 2.275 0.930 ;
        RECT  2.105 1.815 2.275 1.975 ;
        RECT  1.945 1.815 2.105 2.090 ;
        RECT  1.935 1.125 2.095 1.635 ;
        RECT  1.795 0.315 2.055 0.590 ;
        RECT  1.205 1.930 1.945 2.090 ;
        RECT  1.700 1.475 1.935 1.635 ;
        RECT  1.540 1.475 1.700 1.750 ;
        RECT  1.455 0.540 1.615 0.930 ;
        RECT  0.385 1.590 1.540 1.750 ;
        RECT  1.235 0.540 1.455 0.700 ;
        RECT  0.305 0.550 0.385 0.710 ;
        RECT  0.305 1.590 0.385 1.895 ;
        RECT  0.125 0.550 0.305 1.895 ;
    END
END CLKMX2X8MTH

MACRO CLKNAND2X12MTH
    CLASS CORE ;
    FOREIGN CLKNAND2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.965 0.635 5.205 2.100 ;
        RECT  4.570 0.635 4.965 0.935 ;
        RECT  4.685 1.835 4.965 2.100 ;
        RECT  4.385 1.835 4.685 2.505 ;
        RECT  4.270 0.430 4.570 0.935 ;
        RECT  3.725 1.835 4.385 2.425 ;
        RECT  2.075 0.430 4.270 0.730 ;
        RECT  3.465 1.835 3.725 2.485 ;
        RECT  2.805 1.835 3.465 2.425 ;
        RECT  2.505 1.835 2.805 2.505 ;
        RECT  1.875 1.835 2.505 2.425 ;
        RECT  1.575 1.835 1.875 2.505 ;
        RECT  0.965 1.835 1.575 2.425 ;
        RECT  0.665 1.535 0.965 2.425 ;
        RECT  0.265 1.535 0.665 2.235 ;
        END
        AntennaDiffArea 2.241 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.625 1.115 4.785 1.615 ;
        RECT  3.355 1.455 4.625 1.615 ;
        RECT  2.715 1.290 3.355 1.615 ;
        RECT  1.515 1.455 2.715 1.615 ;
        RECT  1.355 1.215 1.515 1.615 ;
        RECT  1.255 1.215 1.355 1.475 ;
        END
        AntennaGateArea 0.8515 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.040 1.115 4.345 1.275 ;
        RECT  3.745 0.920 4.040 1.275 ;
        RECT  2.505 0.950 3.745 1.110 ;
        RECT  1.895 0.950 2.505 1.275 ;
        RECT  1.695 0.875 1.895 1.275 ;
        RECT  0.755 0.875 1.695 1.035 ;
        RECT  0.595 0.875 0.755 1.315 ;
        RECT  0.495 1.055 0.595 1.315 ;
        END
        AntennaGateArea 0.8515 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.070 -0.130 5.330 0.130 ;
        RECT  4.810 -0.130 5.070 0.365 ;
        RECT  3.200 -0.130 4.810 0.130 ;
        RECT  2.940 -0.130 3.200 0.250 ;
        RECT  1.825 -0.130 2.940 0.130 ;
        RECT  1.225 -0.130 1.825 0.640 ;
        RECT  0.725 -0.130 1.225 0.130 ;
        RECT  0.125 -0.130 0.725 0.640 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 2.740 5.330 3.000 ;
        RECT  4.945 2.280 5.205 3.000 ;
        RECT  0.385 2.740 4.945 3.000 ;
        RECT  0.125 2.415 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKNAND2X12MTH

MACRO CLKNAND2X16MTH
    CLASS CORE ;
    FOREIGN CLKNAND2X16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.370 0.430 8.070 2.380 ;
        RECT  1.285 0.430 7.370 0.710 ;
        RECT  7.275 1.495 7.370 2.380 ;
        RECT  4.475 1.760 7.275 2.380 ;
        RECT  3.715 1.760 4.475 2.100 ;
        RECT  3.455 1.760 3.715 2.380 ;
        RECT  2.785 1.760 3.455 2.100 ;
        RECT  2.525 1.760 2.785 2.380 ;
        RECT  1.855 1.760 2.525 2.100 ;
        RECT  1.595 1.760 1.855 2.380 ;
        RECT  0.925 1.760 1.595 2.100 ;
        RECT  0.665 1.760 0.925 2.380 ;
        END
        AntennaDiffArea 3.412 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.055 0.940 7.165 1.100 ;
        RECT  6.895 0.940 7.055 1.540 ;
        RECT  6.145 1.380 6.895 1.540 ;
        RECT  5.545 1.340 6.145 1.540 ;
        RECT  4.395 1.380 5.545 1.540 ;
        RECT  3.750 1.330 4.395 1.540 ;
        RECT  2.570 1.380 3.750 1.540 ;
        RECT  1.970 1.350 2.570 1.540 ;
        RECT  0.755 1.380 1.970 1.540 ;
        RECT  0.495 1.280 0.755 1.540 ;
        END
        AntennaGateArea 1.2896 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.425 0.920 6.685 1.175 ;
        RECT  5.235 0.920 6.425 1.130 ;
        RECT  4.615 0.920 5.235 1.175 ;
        RECT  3.415 0.920 4.615 1.130 ;
        RECT  2.815 0.920 3.415 1.175 ;
        RECT  1.710 0.920 2.815 1.130 ;
        RECT  1.110 0.920 1.710 1.175 ;
        END
        AntennaGateArea 1.2896 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.055 -0.130 8.200 0.130 ;
        RECT  7.115 -0.130 8.055 0.250 ;
        RECT  6.005 -0.130 7.115 0.130 ;
        RECT  5.745 -0.130 6.005 0.250 ;
        RECT  4.145 -0.130 5.745 0.130 ;
        RECT  3.885 -0.130 4.145 0.250 ;
        RECT  2.395 -0.130 3.885 0.130 ;
        RECT  2.135 -0.130 2.395 0.250 ;
        RECT  0.875 -0.130 2.135 0.130 ;
        RECT  0.275 -0.130 0.875 0.690 ;
        RECT  0.000 -0.130 0.275 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 2.740 8.200 3.000 ;
        RECT  7.815 2.570 8.075 3.000 ;
        RECT  4.225 2.740 7.815 3.000 ;
        RECT  3.965 2.300 4.225 3.000 ;
        RECT  0.385 2.740 3.965 3.000 ;
        RECT  0.125 1.820 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKNAND2X16MTH

MACRO CLKNAND2X2MTH
    CLASS CORE ;
    FOREIGN CLKNAND2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.490 0.880 1.540 1.170 ;
        RECT  1.330 0.880 1.490 1.975 ;
        RECT  0.415 0.880 1.330 1.040 ;
        RECT  0.925 1.815 1.330 1.975 ;
        RECT  0.665 1.815 0.925 2.415 ;
        RECT  0.155 0.760 0.415 1.040 ;
        END
        AntennaDiffArea 0.46 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.740 1.245 1.150 1.630 ;
        END
        AntennaGateArea 0.1612 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.450 1.300 0.535 1.560 ;
        RECT  0.180 1.300 0.450 1.990 ;
        RECT  0.100 1.635 0.180 1.990 ;
        END
        AntennaGateArea 0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 -0.130 1.640 0.130 ;
        RECT  1.010 -0.130 1.270 0.690 ;
        RECT  0.760 -0.130 1.010 0.130 ;
        RECT  0.160 -0.130 0.760 0.300 ;
        RECT  0.000 -0.130 0.160 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.470 2.740 1.640 3.000 ;
        RECT  1.210 2.200 1.470 3.000 ;
        RECT  0.385 2.740 1.210 3.000 ;
        RECT  0.125 2.190 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKNAND2X2MTH

MACRO CLKNAND2X4MTH
    CLASS CORE ;
    FOREIGN CLKNAND2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.280 1.290 2.360 1.580 ;
        RECT  2.100 0.515 2.280 2.095 ;
        RECT  1.055 0.515 2.100 0.695 ;
        RECT  1.825 1.915 2.100 2.095 ;
        RECT  1.565 1.915 1.825 2.515 ;
        RECT  0.895 1.915 1.565 2.095 ;
        RECT  0.635 1.915 0.895 2.515 ;
        END
        AntennaDiffArea 0.901 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.755 1.240 1.915 1.735 ;
        RECT  0.775 1.575 1.755 1.735 ;
        RECT  0.460 1.245 0.775 1.735 ;
        END
        AntennaGateArea 0.3185 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 0.880 1.540 1.395 ;
        END
        AntennaGateArea 0.3185 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.165 -0.130 2.460 0.130 ;
        RECT  1.905 -0.130 2.165 0.335 ;
        RECT  0.805 -0.130 1.905 0.130 ;
        RECT  0.205 -0.130 0.805 0.685 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  2.075 2.295 2.335 3.000 ;
        RECT  0.385 2.740 2.075 3.000 ;
        RECT  0.125 1.925 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKNAND2X4MTH

MACRO CLKNAND2X8MTH
    CLASS CORE ;
    FOREIGN CLKNAND2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.315 1.495 4.410 2.315 ;
        RECT  4.045 0.430 4.315 2.315 ;
        RECT  1.125 0.430 4.045 0.700 ;
        RECT  3.845 1.965 4.045 2.315 ;
        RECT  3.585 1.965 3.845 2.465 ;
        RECT  2.875 1.965 3.585 2.315 ;
        RECT  2.615 1.965 2.875 2.465 ;
        RECT  1.895 1.965 2.615 2.315 ;
        RECT  1.635 1.965 1.895 2.465 ;
        RECT  0.925 1.965 1.635 2.315 ;
        RECT  0.665 1.965 0.925 2.465 ;
        END
        AntennaDiffArea 1.683 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.645 1.025 3.865 1.745 ;
        RECT  2.555 1.585 3.645 1.745 ;
        RECT  1.915 1.265 2.555 1.745 ;
        RECT  0.685 1.585 1.915 1.745 ;
        RECT  0.525 1.255 0.685 1.745 ;
        RECT  0.425 1.255 0.525 1.515 ;
        END
        AntennaGateArea 0.6396 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.145 3.370 1.405 ;
        RECT  2.770 0.920 3.220 1.405 ;
        RECT  1.555 0.920 2.770 1.080 ;
        RECT  1.395 0.920 1.555 1.385 ;
        RECT  1.295 1.125 1.395 1.385 ;
        END
        AntennaGateArea 0.6396 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.115 -0.130 4.510 0.130 ;
        RECT  3.855 -0.130 4.115 0.250 ;
        RECT  2.285 -0.130 3.855 0.130 ;
        RECT  2.025 -0.130 2.285 0.250 ;
        RECT  0.805 -0.130 2.025 0.130 ;
        RECT  0.205 -0.130 0.805 0.690 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 2.540 4.385 3.000 ;
        RECT  0.385 2.740 4.125 3.000 ;
        RECT  0.125 1.925 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END CLKNAND2X8MTH

MACRO CLKXOR2X12MTH
    CLASS CORE ;
    FOREIGN CLKXOR2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.325 1.125 12.585 2.385 ;
        RECT  11.505 1.125 12.325 1.955 ;
        RECT  11.495 1.125 11.505 2.450 ;
        RECT  11.245 0.435 11.495 2.450 ;
        RECT  11.005 0.435 11.245 2.125 ;
        RECT  9.955 0.435 11.005 0.925 ;
        RECT  10.575 1.525 11.005 2.125 ;
        RECT  10.315 1.525 10.575 2.490 ;
        END
        AntennaDiffArea 1.48 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.615 1.290 2.370 1.550 ;
        END
        AntennaGateArea 0.7644 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.625 0.900 9.575 1.195 ;
        END
        AntennaGateArea 0.7631 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.275 -0.130 12.710 0.130 ;
        RECT  11.675 -0.130 12.275 0.665 ;
        RECT  10.855 -0.130 11.675 0.130 ;
        RECT  10.595 -0.130 10.855 0.250 ;
        RECT  9.775 -0.130 10.595 0.130 ;
        RECT  9.175 -0.130 9.775 0.690 ;
        RECT  3.850 -0.130 9.175 0.130 ;
        RECT  3.590 -0.130 3.850 0.785 ;
        RECT  2.770 -0.130 3.590 0.130 ;
        RECT  2.510 -0.130 2.770 0.765 ;
        RECT  2.005 -0.130 2.510 0.130 ;
        RECT  1.745 -0.130 2.005 0.765 ;
        RECT  0.925 -0.130 1.745 0.130 ;
        RECT  0.665 -0.130 0.925 0.765 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.045 2.740 12.710 3.000 ;
        RECT  11.785 2.135 12.045 3.000 ;
        RECT  10.035 2.740 11.785 3.000 ;
        RECT  9.775 2.570 10.035 3.000 ;
        RECT  1.915 2.740 9.775 3.000 ;
        RECT  1.655 2.085 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.105 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.045 1.135 10.825 1.295 ;
        RECT  9.885 1.135 10.045 2.180 ;
        RECT  8.985 2.020 9.885 2.180 ;
        RECT  9.395 1.570 9.495 1.830 ;
        RECT  9.235 1.380 9.395 1.830 ;
        RECT  8.445 1.380 9.235 1.540 ;
        RECT  8.725 1.735 8.985 2.335 ;
        RECT  8.445 0.460 8.895 0.720 ;
        RECT  7.970 1.735 8.725 1.895 ;
        RECT  8.215 2.200 8.475 2.560 ;
        RECT  8.185 0.460 8.445 1.540 ;
        RECT  7.455 2.400 8.215 2.560 ;
        RECT  7.810 0.310 7.970 2.035 ;
        RECT  7.090 0.310 7.810 0.470 ;
        RECT  7.785 1.735 7.810 2.035 ;
        RECT  7.705 1.775 7.785 2.035 ;
        RECT  7.455 0.655 7.630 0.915 ;
        RECT  7.295 0.655 7.455 2.560 ;
        RECT  6.550 1.095 7.295 1.255 ;
        RECT  7.195 1.835 7.295 2.560 ;
        RECT  2.895 2.400 7.195 2.560 ;
        RECT  6.830 0.310 7.090 0.915 ;
        RECT  6.845 1.835 6.945 2.095 ;
        RECT  6.685 1.620 6.845 2.095 ;
        RECT  6.040 0.310 6.830 0.470 ;
        RECT  5.940 1.620 6.685 1.780 ;
        RECT  6.390 0.735 6.550 1.255 ;
        RECT  6.175 1.960 6.435 2.220 ;
        RECT  6.290 0.735 6.390 0.995 ;
        RECT  5.355 2.060 6.175 2.220 ;
        RECT  5.940 0.310 6.040 0.950 ;
        RECT  5.780 0.310 5.940 1.880 ;
        RECT  4.930 0.310 5.780 0.470 ;
        RECT  5.635 1.575 5.780 1.880 ;
        RECT  5.355 0.655 5.470 0.915 ;
        RECT  5.195 0.655 5.355 2.220 ;
        RECT  5.095 1.960 5.195 2.220 ;
        RECT  4.335 2.060 5.095 2.220 ;
        RECT  4.770 0.310 4.930 0.805 ;
        RECT  4.770 1.720 4.815 1.880 ;
        RECT  4.610 0.545 4.770 1.880 ;
        RECT  4.555 1.720 4.610 1.880 ;
        RECT  4.335 0.525 4.390 0.785 ;
        RECT  4.175 0.525 4.335 2.220 ;
        RECT  4.130 0.525 4.175 0.785 ;
        RECT  4.045 1.620 4.175 2.220 ;
        RECT  3.365 2.060 4.045 2.220 ;
        RECT  3.205 0.525 3.365 2.220 ;
        RECT  3.050 0.525 3.205 0.785 ;
        RECT  3.105 1.620 3.205 2.220 ;
        RECT  2.895 1.010 3.025 1.270 ;
        RECT  2.735 0.945 2.895 2.560 ;
        RECT  1.465 0.945 2.735 1.105 ;
        RECT  2.425 1.730 2.735 1.890 ;
        RECT  2.165 1.730 2.425 2.330 ;
        RECT  1.405 1.730 2.165 1.890 ;
        RECT  1.205 0.715 1.465 1.105 ;
        RECT  1.145 1.730 1.405 2.330 ;
        RECT  0.385 0.945 1.205 1.105 ;
        RECT  0.385 1.730 1.145 1.890 ;
        RECT  0.125 0.715 0.385 1.105 ;
        RECT  0.125 1.730 0.385 2.330 ;
    END
END CLKXOR2X12MTH

MACRO CLKXOR2X16MTH
    CLASS CORE ;
    FOREIGN CLKXOR2X16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.990 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.605 0.520 15.865 2.385 ;
        RECT  14.785 1.085 15.605 1.785 ;
        RECT  14.745 1.085 14.785 2.385 ;
        RECT  14.525 0.470 14.745 2.385 ;
        RECT  14.485 0.470 14.525 1.785 ;
        RECT  13.825 1.085 14.485 1.785 ;
        RECT  13.665 1.085 13.825 2.385 ;
        RECT  13.565 0.495 13.665 2.385 ;
        RECT  13.405 0.495 13.565 2.045 ;
        RECT  12.885 1.785 13.405 2.045 ;
        RECT  12.625 1.785 12.885 2.385 ;
        END
        AntennaDiffArea 1.999 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.515 1.285 3.055 1.550 ;
        END
        AntennaGateArea 1.0205 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.710 1.045 11.310 1.540 ;
        RECT  10.415 1.045 10.710 1.205 ;
        END
        AntennaGateArea 1.0101 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.285 -0.130 15.990 0.130 ;
        RECT  15.025 -0.130 15.285 0.805 ;
        RECT  14.205 -0.130 15.025 0.130 ;
        RECT  13.945 -0.130 14.205 0.815 ;
        RECT  13.125 -0.130 13.945 0.130 ;
        RECT  12.865 -0.130 13.125 0.675 ;
        RECT  12.585 -0.130 12.865 0.130 ;
        RECT  12.325 -0.130 12.585 0.520 ;
        RECT  11.445 -0.130 12.325 0.130 ;
        RECT  11.185 -0.130 11.445 0.515 ;
        RECT  5.570 -0.130 11.185 0.130 ;
        RECT  5.310 -0.130 5.570 0.300 ;
        RECT  4.440 -0.130 5.310 0.130 ;
        RECT  4.180 -0.130 4.440 0.300 ;
        RECT  3.360 -0.130 4.180 0.130 ;
        RECT  3.100 -0.130 3.360 0.765 ;
        RECT  2.825 -0.130 3.100 0.130 ;
        RECT  2.565 -0.130 2.825 0.765 ;
        RECT  1.745 -0.130 2.565 0.130 ;
        RECT  1.485 -0.130 1.745 0.765 ;
        RECT  0.665 -0.130 1.485 0.130 ;
        RECT  0.405 -0.130 0.665 0.990 ;
        RECT  0.000 -0.130 0.405 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.325 2.740 15.990 3.000 ;
        RECT  15.065 2.120 15.325 3.000 ;
        RECT  12.345 2.740 15.065 3.000 ;
        RECT  12.085 2.220 12.345 3.000 ;
        RECT  2.775 2.740 12.085 3.000 ;
        RECT  2.515 2.085 2.775 3.000 ;
        RECT  0.000 2.740 2.515 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.365 1.120 13.165 1.380 ;
        RECT  12.205 1.120 12.365 2.015 ;
        RECT  10.785 1.855 12.205 2.015 ;
        RECT  11.805 0.355 12.015 0.855 ;
        RECT  11.755 0.355 11.805 1.670 ;
        RECT  11.545 0.695 11.755 1.670 ;
        RECT  10.875 0.695 11.545 0.855 ;
        RECT  11.035 2.200 11.295 2.560 ;
        RECT  10.275 2.400 11.035 2.560 ;
        RECT  10.615 0.355 10.875 0.855 ;
        RECT  10.525 1.775 10.785 2.165 ;
        RECT  10.175 0.695 10.615 0.855 ;
        RECT  9.765 1.775 10.525 1.935 ;
        RECT  10.015 2.200 10.275 2.560 ;
        RECT  9.955 0.695 10.175 1.170 ;
        RECT  9.255 2.400 10.015 2.560 ;
        RECT  9.665 0.655 9.775 0.915 ;
        RECT  9.665 1.775 9.765 2.035 ;
        RECT  9.505 0.310 9.665 2.035 ;
        RECT  8.805 0.310 9.505 0.470 ;
        RECT  9.255 0.655 9.315 0.915 ;
        RECT  8.995 0.655 9.255 2.560 ;
        RECT  8.295 1.095 8.995 1.255 ;
        RECT  3.435 2.400 8.995 2.560 ;
        RECT  8.545 0.310 8.805 0.915 ;
        RECT  8.645 1.835 8.745 2.095 ;
        RECT  8.485 1.620 8.645 2.095 ;
        RECT  7.785 0.310 8.545 0.470 ;
        RECT  7.740 1.620 8.485 1.780 ;
        RECT  8.135 0.735 8.295 1.255 ;
        RECT  7.975 1.960 8.235 2.220 ;
        RECT  8.035 0.735 8.135 0.995 ;
        RECT  7.155 2.060 7.975 2.220 ;
        RECT  7.595 0.310 7.785 0.950 ;
        RECT  7.595 1.620 7.740 1.880 ;
        RECT  7.435 0.310 7.595 1.880 ;
        RECT  6.695 0.310 7.435 0.470 ;
        RECT  7.105 0.650 7.245 0.810 ;
        RECT  7.105 1.960 7.155 2.220 ;
        RECT  6.945 0.650 7.105 2.220 ;
        RECT  6.895 1.960 6.945 2.220 ;
        RECT  6.075 2.060 6.895 2.220 ;
        RECT  6.615 0.310 6.695 0.805 ;
        RECT  6.455 0.310 6.615 1.880 ;
        RECT  6.355 1.720 6.455 1.880 ;
        RECT  5.165 0.525 6.225 0.785 ;
        RECT  5.815 1.960 6.075 2.220 ;
        RECT  5.165 2.060 5.815 2.220 ;
        RECT  4.905 0.525 5.165 2.220 ;
        RECT  3.640 0.525 4.905 0.785 ;
        RECT  4.225 2.060 4.905 2.220 ;
        RECT  3.435 1.010 4.615 1.270 ;
        RECT  3.965 1.620 4.225 2.220 ;
        RECT  3.275 0.945 3.435 2.560 ;
        RECT  2.285 0.945 3.275 1.105 ;
        RECT  3.025 1.730 3.275 2.330 ;
        RECT  2.265 1.730 3.025 1.890 ;
        RECT  2.025 0.715 2.285 1.105 ;
        RECT  2.005 1.730 2.265 2.330 ;
        RECT  1.205 0.945 2.025 1.105 ;
        RECT  1.325 1.730 2.005 1.890 ;
        RECT  1.065 1.730 1.325 2.330 ;
        RECT  0.945 0.715 1.205 1.105 ;
        RECT  0.385 1.730 1.065 1.890 ;
        RECT  0.125 1.730 0.385 2.330 ;
    END
END CLKXOR2X16MTH

MACRO CLKXOR2X2MTH
    CLASS CORE ;
    FOREIGN CLKXOR2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.845 0.470 4.005 2.425 ;
        RECT  3.715 0.470 3.845 1.025 ;
        RECT  3.715 2.165 3.845 2.425 ;
        END
        AntennaDiffArea 0.401 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.585 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 1.185 3.270 1.580 ;
        END
        AntennaGateArea 0.1859 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.825 -0.130 4.100 0.130 ;
        RECT  3.225 -0.130 3.825 0.290 ;
        RECT  0.615 -0.130 3.225 0.130 ;
        RECT  0.355 -0.130 0.615 0.300 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  2.835 2.620 3.435 3.000 ;
        RECT  1.605 2.740 2.835 3.000 ;
        RECT  0.665 2.570 1.605 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.505 1.215 3.665 1.975 ;
        RECT  3.355 1.815 3.505 1.975 ;
        RECT  3.195 1.815 3.355 2.405 ;
        RECT  2.680 2.245 3.195 2.405 ;
        RECT  2.755 1.800 2.945 2.060 ;
        RECT  2.755 0.765 2.845 1.025 ;
        RECT  2.595 0.765 2.755 2.060 ;
        RECT  2.520 2.245 2.680 2.455 ;
        RECT  2.545 1.270 2.595 1.530 ;
        RECT  1.925 2.295 2.520 2.455 ;
        RECT  2.335 0.365 2.385 0.625 ;
        RECT  2.335 1.855 2.385 2.115 ;
        RECT  2.175 0.365 2.335 2.115 ;
        RECT  2.125 0.365 2.175 0.625 ;
        RECT  0.945 0.365 2.125 0.525 ;
        RECT  1.925 0.830 1.955 1.090 ;
        RECT  1.765 0.830 1.925 2.455 ;
        RECT  1.695 0.830 1.765 1.090 ;
        RECT  1.665 1.980 1.765 2.240 ;
        RECT  1.195 0.765 1.355 2.145 ;
        RECT  1.135 0.765 1.195 1.025 ;
        RECT  0.945 1.225 1.015 1.485 ;
        RECT  0.785 0.365 0.945 1.920 ;
        RECT  0.385 0.865 0.785 1.025 ;
        RECT  0.385 1.760 0.785 1.920 ;
        RECT  0.125 0.765 0.385 1.025 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END CLKXOR2X2MTH

MACRO CLKXOR2X4MTH
    CLASS CORE ;
    FOREIGN CLKXOR2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.995 0.580 6.165 0.840 ;
        RECT  5.995 1.290 6.050 1.580 ;
        RECT  5.815 0.580 5.995 2.385 ;
        RECT  5.665 1.785 5.815 2.385 ;
        END
        AntennaDiffArea 0.541 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.220 0.955 1.550 ;
        RECT  0.100 1.220 0.310 1.580 ;
        END
        AntennaGateArea 0.2535 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.375 1.110 4.535 1.370 ;
        RECT  3.930 1.210 4.375 1.370 ;
        RECT  3.770 1.210 3.930 2.220 ;
        RECT  3.545 1.210 3.770 1.370 ;
        RECT  2.225 2.060 3.770 2.220 ;
        RECT  3.545 0.310 3.590 0.470 ;
        RECT  3.385 0.310 3.545 1.370 ;
        RECT  3.330 0.310 3.385 0.470 ;
        RECT  2.225 1.205 2.400 1.540 ;
        RECT  2.065 1.205 2.225 2.220 ;
        RECT  1.905 1.205 2.065 1.540 ;
        END
        AntennaGateArea 0.2834 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.635 -0.130 6.560 0.130 ;
        RECT  5.395 -0.130 5.635 0.820 ;
        RECT  5.025 -0.130 5.395 0.250 ;
        RECT  4.710 -0.130 5.025 0.130 ;
        RECT  3.770 -0.130 4.710 0.250 ;
        RECT  2.955 -0.130 3.770 0.130 ;
        RECT  2.015 -0.130 2.955 0.250 ;
        RECT  1.780 -0.130 2.015 0.130 ;
        RECT  1.520 -0.130 1.780 0.250 ;
        RECT  0.705 -0.130 1.520 0.130 ;
        RECT  0.415 -0.130 0.705 0.925 ;
        RECT  0.000 -0.130 0.415 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.785 6.435 3.000 ;
        RECT  1.530 2.740 6.175 3.000 ;
        RECT  1.270 2.570 1.530 3.000 ;
        RECT  0.000 2.740 1.270 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.215 1.220 5.545 1.480 ;
        RECT  5.055 0.430 5.215 2.050 ;
        RECT  3.930 0.430 5.055 0.590 ;
        RECT  5.015 1.890 5.055 2.050 ;
        RECT  4.755 1.890 5.015 2.150 ;
        RECT  4.715 0.770 4.875 1.710 ;
        RECT  4.185 0.770 4.715 0.930 ;
        RECT  4.490 1.550 4.715 1.710 ;
        RECT  4.330 1.550 4.490 2.560 ;
        RECT  4.240 1.890 4.330 2.560 ;
        RECT  1.885 2.400 4.240 2.560 ;
        RECT  3.770 0.430 3.930 0.940 ;
        RECT  3.725 0.680 3.770 0.940 ;
        RECT  3.150 1.720 3.575 1.880 ;
        RECT  3.150 0.660 3.205 0.920 ;
        RECT  2.990 0.430 3.150 1.880 ;
        RECT  1.725 0.430 2.990 0.590 ;
        RECT  2.745 1.230 2.810 1.490 ;
        RECT  2.585 0.770 2.745 1.880 ;
        RECT  2.485 0.770 2.585 0.930 ;
        RECT  2.405 1.720 2.585 1.880 ;
        RECT  1.725 2.170 1.885 2.560 ;
        RECT  1.565 0.430 1.725 1.980 ;
        RECT  1.335 2.170 1.725 2.330 ;
        RECT  1.515 0.700 1.565 0.960 ;
        RECT  1.515 1.720 1.565 1.980 ;
        RECT  1.335 1.225 1.385 1.485 ;
        RECT  1.215 0.815 1.335 2.330 ;
        RECT  1.175 0.715 1.215 2.330 ;
        RECT  0.955 0.715 1.175 0.975 ;
        RECT  0.525 1.730 1.175 2.330 ;
    END
END CLKXOR2X4MTH

MACRO CLKXOR2X8MTH
    CLASS CORE ;
    FOREIGN CLKXOR2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.945 1.260 9.205 2.385 ;
        RECT  8.185 1.260 8.945 1.610 ;
        RECT  7.920 0.625 8.185 2.385 ;
        END
        AntennaDiffArea 0.906 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.275 1.745 1.545 ;
        END
        AntennaGateArea 0.507 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.310 1.015 3.370 1.275 ;
        RECT  2.970 1.015 3.310 1.580 ;
        END
        AntennaGateArea 0.507 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.060 -0.130 9.840 0.130 ;
        RECT  8.460 -0.130 9.060 0.980 ;
        RECT  7.640 -0.130 8.460 0.130 ;
        RECT  7.040 -0.130 7.640 0.980 ;
        RECT  3.135 -0.130 7.040 0.130 ;
        RECT  2.875 -0.130 3.135 0.740 ;
        RECT  1.990 -0.130 2.875 0.130 ;
        RECT  1.390 -0.130 1.990 0.690 ;
        RECT  0.510 -0.130 1.390 0.130 ;
        RECT  0.250 -0.130 0.510 0.990 ;
        RECT  0.000 -0.130 0.250 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.715 2.740 9.840 3.000 ;
        RECT  9.455 1.905 9.715 3.000 ;
        RECT  8.695 2.740 9.455 3.000 ;
        RECT  8.435 1.835 8.695 3.000 ;
        RECT  7.645 2.740 8.435 3.000 ;
        RECT  7.385 2.570 7.645 3.000 ;
        RECT  0.385 2.740 7.385 3.000 ;
        RECT  0.125 1.765 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.430 1.220 7.690 1.480 ;
        RECT  6.715 1.320 7.430 1.480 ;
        RECT  7.175 1.700 7.275 2.300 ;
        RECT  7.015 1.700 7.175 2.540 ;
        RECT  6.255 2.380 7.015 2.540 ;
        RECT  6.715 1.840 6.765 2.100 ;
        RECT  6.555 0.560 6.715 2.100 ;
        RECT  6.410 0.560 6.555 0.720 ;
        RECT  6.505 1.840 6.555 2.100 ;
        RECT  6.150 0.310 6.410 0.720 ;
        RECT  6.155 2.010 6.255 2.540 ;
        RECT  5.995 0.900 6.155 2.540 ;
        RECT  5.300 0.310 6.150 0.470 ;
        RECT  5.870 0.900 5.995 1.060 ;
        RECT  2.220 2.380 5.995 2.540 ;
        RECT  5.710 0.650 5.870 1.060 ;
        RECT  5.485 1.665 5.745 1.860 ;
        RECT  5.610 0.650 5.710 0.810 ;
        RECT  5.300 1.665 5.485 1.825 ;
        RECT  5.140 0.310 5.300 1.825 ;
        RECT  4.975 2.005 5.235 2.200 ;
        RECT  5.040 0.310 5.140 0.740 ;
        RECT  4.465 1.665 5.140 1.825 ;
        RECT  4.220 0.310 5.040 0.470 ;
        RECT  4.220 2.040 4.975 2.200 ;
        RECT  4.635 0.650 4.760 0.810 ;
        RECT  4.475 0.650 4.635 1.375 ;
        RECT  4.220 1.215 4.475 1.375 ;
        RECT  4.060 0.310 4.220 0.745 ;
        RECT  4.060 1.215 4.220 2.200 ;
        RECT  3.960 0.485 4.060 0.745 ;
        RECT  3.955 1.600 4.060 2.200 ;
        RECT  2.765 2.040 3.955 2.200 ;
        RECT  3.710 1.140 3.880 1.400 ;
        RECT  3.550 0.535 3.710 1.860 ;
        RECT  3.445 0.535 3.550 0.795 ;
        RECT  3.445 1.700 3.550 1.860 ;
        RECT  2.660 1.575 2.765 2.200 ;
        RECT  2.500 0.470 2.660 2.200 ;
        RECT  2.335 0.470 2.500 0.730 ;
        RECT  2.220 0.925 2.320 1.185 ;
        RECT  2.060 0.925 2.220 2.540 ;
        RECT  1.050 0.925 2.060 1.085 ;
        RECT  0.635 1.765 2.060 2.365 ;
        RECT  0.790 0.715 1.050 1.085 ;
    END
END CLKXOR2X8MTH

MACRO DFFHQNX1MTH
    CLASS CORE ;
    FOREIGN DFFHQNX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.735 8.920 2.125 ;
        RECT  8.635 0.735 8.710 0.995 ;
        RECT  8.635 1.865 8.710 2.125 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 0.880 2.360 1.445 ;
        RECT  2.030 1.185 2.105 1.445 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.145 0.765 1.595 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.805 -0.130 9.020 0.130 ;
        RECT  8.305 -0.130 8.805 0.415 ;
        RECT  7.565 -0.130 8.305 0.130 ;
        RECT  7.305 -0.130 7.565 0.250 ;
        RECT  6.150 -0.130 7.305 0.130 ;
        RECT  5.550 -0.130 6.150 0.250 ;
        RECT  4.680 -0.130 5.550 0.130 ;
        RECT  3.740 -0.130 4.680 0.250 ;
        RECT  2.430 -0.130 3.740 0.130 ;
        RECT  2.270 -0.130 2.430 0.700 ;
        RECT  0.530 -0.130 2.270 0.130 ;
        RECT  0.270 -0.130 0.530 0.250 ;
        RECT  0.000 -0.130 0.270 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.865 2.740 9.020 3.000 ;
        RECT  8.265 2.620 8.865 3.000 ;
        RECT  5.855 2.740 8.265 3.000 ;
        RECT  4.915 2.620 5.855 3.000 ;
        RECT  0.765 2.740 4.915 3.000 ;
        RECT  0.165 2.405 0.765 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.875 1.290 8.460 1.550 ;
        RECT  7.475 0.430 8.125 0.590 ;
        RECT  7.535 2.320 8.125 2.480 ;
        RECT  7.875 0.800 7.925 0.960 ;
        RECT  7.715 0.800 7.875 2.140 ;
        RECT  7.665 0.800 7.715 0.960 ;
        RECT  7.475 1.210 7.535 2.480 ;
        RECT  7.375 0.430 7.475 2.480 ;
        RECT  7.315 0.430 7.375 1.370 ;
        RECT  6.845 2.000 7.375 2.210 ;
        RECT  7.030 0.430 7.315 0.590 ;
        RECT  7.035 1.520 7.195 1.780 ;
        RECT  6.735 1.520 7.035 1.680 ;
        RECT  6.770 0.355 7.030 0.590 ;
        RECT  6.685 1.950 6.845 2.210 ;
        RECT  6.585 1.475 6.735 1.680 ;
        RECT  6.575 0.430 6.585 1.680 ;
        RECT  6.425 0.430 6.575 1.635 ;
        RECT  6.505 2.370 6.555 2.530 ;
        RECT  6.295 2.280 6.505 2.530 ;
        RECT  5.120 0.430 6.425 0.590 ;
        RECT  5.985 1.475 6.425 1.635 ;
        RECT  4.645 2.280 6.295 2.440 ;
        RECT  5.805 1.940 6.285 2.100 ;
        RECT  5.805 0.785 6.240 0.945 ;
        RECT  5.645 0.785 5.805 2.100 ;
        RECT  4.985 1.940 5.645 2.100 ;
        RECT  5.325 1.570 5.465 1.730 ;
        RECT  5.165 0.770 5.325 1.730 ;
        RECT  4.095 0.770 5.165 0.930 ;
        RECT  4.860 0.350 5.120 0.590 ;
        RECT  4.825 1.280 4.985 2.100 ;
        RECT  3.740 0.430 4.860 0.590 ;
        RECT  4.705 1.280 4.825 1.440 ;
        RECT  4.485 1.650 4.645 2.540 ;
        RECT  4.435 1.650 4.485 1.810 ;
        RECT  3.800 2.380 4.485 2.540 ;
        RECT  4.275 1.550 4.435 1.810 ;
        RECT  4.095 1.990 4.285 2.150 ;
        RECT  3.935 0.770 4.095 2.150 ;
        RECT  3.410 0.990 3.935 1.190 ;
        RECT  3.640 2.355 3.800 2.540 ;
        RECT  3.580 0.430 3.740 0.810 ;
        RECT  1.105 2.355 3.640 2.515 ;
        RECT  3.110 0.650 3.580 0.810 ;
        RECT  2.770 0.310 3.400 0.470 ;
        RECT  3.110 1.255 3.220 1.515 ;
        RECT  2.950 0.650 3.110 2.175 ;
        RECT  1.445 2.015 2.950 2.175 ;
        RECT  2.610 0.310 2.770 1.835 ;
        RECT  1.850 1.675 2.610 1.835 ;
        RECT  1.850 0.755 1.895 0.915 ;
        RECT  1.690 0.755 1.850 1.835 ;
        RECT  1.525 0.385 1.785 0.575 ;
        RECT  1.635 0.755 1.690 0.915 ;
        RECT  0.765 0.415 1.525 0.575 ;
        RECT  1.285 1.395 1.445 2.175 ;
        RECT  1.105 0.755 1.385 0.915 ;
        RECT  0.945 0.755 1.105 2.515 ;
        RECT  0.605 0.415 0.765 0.865 ;
        RECT  0.385 0.705 0.605 0.865 ;
        RECT  0.285 0.705 0.385 0.965 ;
        RECT  0.285 1.795 0.385 2.055 ;
        RECT  0.125 0.705 0.285 2.055 ;
    END
END DFFHQNX1MTH

MACRO DFFHQNX2MTH
    CLASS CORE ;
    FOREIGN DFFHQNX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 2.080 8.920 2.400 ;
        RECT  8.735 0.425 8.895 2.400 ;
        RECT  8.635 0.425 8.735 1.025 ;
        RECT  8.635 1.785 8.735 2.400 ;
        END
        AntennaDiffArea 0.521 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 0.880 2.445 1.445 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.130 0.765 1.580 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.345 -0.130 9.020 0.130 ;
        RECT  8.085 -0.130 8.345 0.250 ;
        RECT  7.565 -0.130 8.085 0.130 ;
        RECT  7.305 -0.130 7.565 0.250 ;
        RECT  6.265 -0.130 7.305 0.130 ;
        RECT  5.325 -0.130 6.265 0.250 ;
        RECT  4.560 -0.130 5.325 0.130 ;
        RECT  3.620 -0.130 4.560 0.250 ;
        RECT  2.445 -0.130 3.620 0.130 ;
        RECT  2.285 -0.130 2.445 0.700 ;
        RECT  0.605 -0.130 2.285 0.130 ;
        RECT  0.345 -0.130 0.605 0.250 ;
        RECT  0.000 -0.130 0.345 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.275 2.740 9.020 3.000 ;
        RECT  7.675 2.580 8.275 3.000 ;
        RECT  5.855 2.740 7.675 3.000 ;
        RECT  4.915 2.620 5.855 3.000 ;
        RECT  0.945 2.740 4.915 3.000 ;
        RECT  0.345 2.365 0.945 3.000 ;
        RECT  0.000 2.740 0.345 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.875 1.255 8.555 1.515 ;
        RECT  7.535 2.240 8.095 2.400 ;
        RECT  7.875 0.770 7.925 0.930 ;
        RECT  7.745 0.310 7.905 0.590 ;
        RECT  7.715 0.770 7.875 2.060 ;
        RECT  7.475 0.430 7.745 0.590 ;
        RECT  7.665 0.770 7.715 0.930 ;
        RECT  7.475 1.210 7.535 2.400 ;
        RECT  7.375 0.430 7.475 2.400 ;
        RECT  7.315 0.430 7.375 1.370 ;
        RECT  6.685 1.950 7.375 2.210 ;
        RECT  7.030 0.430 7.315 0.590 ;
        RECT  7.035 1.510 7.195 1.770 ;
        RECT  6.585 1.510 7.035 1.670 ;
        RECT  6.770 0.355 7.030 0.590 ;
        RECT  6.425 0.430 6.585 1.670 ;
        RECT  6.455 2.370 6.555 2.530 ;
        RECT  6.295 2.280 6.455 2.530 ;
        RECT  5.135 0.430 6.425 0.590 ;
        RECT  5.985 1.470 6.425 1.670 ;
        RECT  5.805 1.940 6.295 2.100 ;
        RECT  4.650 2.280 6.295 2.440 ;
        RECT  5.805 0.785 6.245 0.945 ;
        RECT  5.645 0.785 5.805 2.100 ;
        RECT  4.990 1.940 5.645 2.100 ;
        RECT  5.330 1.560 5.465 1.720 ;
        RECT  5.170 0.770 5.330 1.720 ;
        RECT  4.045 0.770 5.170 0.930 ;
        RECT  4.875 0.310 5.135 0.590 ;
        RECT  4.830 1.140 4.990 2.100 ;
        RECT  3.705 0.430 4.875 0.590 ;
        RECT  4.570 1.140 4.830 1.300 ;
        RECT  4.490 1.620 4.650 2.560 ;
        RECT  4.225 1.620 4.490 1.780 ;
        RECT  3.370 2.400 4.490 2.560 ;
        RECT  4.045 2.010 4.285 2.170 ;
        RECT  3.885 0.770 4.045 2.170 ;
        RECT  3.425 0.990 3.885 1.190 ;
        RECT  3.545 0.430 3.705 0.810 ;
        RECT  3.125 0.650 3.545 0.810 ;
        RECT  3.125 1.495 3.525 1.755 ;
        RECT  3.210 2.355 3.370 2.560 ;
        RECT  2.785 0.310 3.365 0.470 ;
        RECT  1.285 2.355 3.210 2.515 ;
        RECT  2.965 0.650 3.125 2.175 ;
        RECT  1.625 2.015 2.965 2.175 ;
        RECT  2.625 0.310 2.785 1.835 ;
        RECT  1.965 1.675 2.625 1.835 ;
        RECT  1.805 0.755 1.965 1.835 ;
        RECT  1.555 0.310 1.815 0.575 ;
        RECT  1.665 0.755 1.805 0.915 ;
        RECT  1.465 1.735 1.625 2.175 ;
        RECT  0.945 0.415 1.555 0.575 ;
        RECT  1.285 0.755 1.415 0.915 ;
        RECT  1.125 0.755 1.285 2.515 ;
        RECT  0.785 0.415 0.945 0.865 ;
        RECT  0.385 0.705 0.785 0.865 ;
        RECT  0.285 0.705 0.385 0.965 ;
        RECT  0.285 1.760 0.385 2.020 ;
        RECT  0.125 0.705 0.285 2.020 ;
    END
END DFFHQNX2MTH

MACRO DFFHQNX4MTH
    CLASS CORE ;
    FOREIGN DFFHQNX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.990 1.700 8.285 2.315 ;
        RECT  7.990 0.770 8.225 0.950 ;
        RECT  7.810 0.770 7.990 2.315 ;
        END
        AntennaDiffArea 0.582 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 0.880 2.360 1.445 ;
        RECT  2.005 1.185 2.105 1.445 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.210 0.765 1.740 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 -0.130 9.430 0.130 ;
        RECT  9.045 -0.130 9.305 0.300 ;
        RECT  7.615 -0.130 9.045 0.130 ;
        RECT  7.355 -0.130 7.615 0.250 ;
        RECT  6.255 -0.130 7.355 0.130 ;
        RECT  5.315 -0.130 6.255 0.250 ;
        RECT  4.570 -0.130 5.315 0.130 ;
        RECT  3.630 -0.130 4.570 0.250 ;
        RECT  2.415 -0.130 3.630 0.130 ;
        RECT  2.215 -0.130 2.415 0.700 ;
        RECT  0.605 -0.130 2.215 0.130 ;
        RECT  0.345 -0.130 0.605 0.250 ;
        RECT  0.000 -0.130 0.345 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.205 2.740 9.430 3.000 ;
        RECT  8.605 2.570 9.205 3.000 ;
        RECT  7.785 2.740 8.605 3.000 ;
        RECT  6.845 2.570 7.785 3.000 ;
        RECT  5.855 2.740 6.845 3.000 ;
        RECT  4.915 2.620 5.855 3.000 ;
        RECT  0.765 2.740 4.915 3.000 ;
        RECT  0.165 2.455 0.765 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.145 0.565 9.305 2.055 ;
        RECT  9.025 0.565 9.145 0.825 ;
        RECT  9.045 1.715 9.145 2.055 ;
        RECT  8.625 1.715 9.045 1.875 ;
        RECT  8.805 1.010 8.965 1.500 ;
        RECT  8.725 1.010 8.805 1.170 ;
        RECT  8.565 0.430 8.725 1.170 ;
        RECT  8.465 1.355 8.625 1.875 ;
        RECT  7.535 0.430 8.565 0.590 ;
        RECT  8.430 1.355 8.465 1.515 ;
        RECT  8.170 1.310 8.430 1.515 ;
        RECT  7.375 0.430 7.535 2.210 ;
        RECT  6.925 0.430 7.375 0.590 ;
        RECT  6.895 2.050 7.375 2.210 ;
        RECT  6.585 1.445 7.195 1.720 ;
        RECT  6.765 0.365 6.925 0.625 ;
        RECT  6.635 1.950 6.895 2.210 ;
        RECT  6.425 0.430 6.585 1.720 ;
        RECT  6.465 2.400 6.555 2.560 ;
        RECT  6.205 2.280 6.465 2.560 ;
        RECT  5.135 0.430 6.425 0.590 ;
        RECT  5.985 1.460 6.425 1.720 ;
        RECT  5.805 0.815 6.245 0.975 ;
        RECT  5.805 1.940 6.210 2.100 ;
        RECT  4.655 2.280 6.205 2.440 ;
        RECT  5.645 0.815 5.805 2.100 ;
        RECT  4.995 1.940 5.645 2.100 ;
        RECT  5.335 1.600 5.465 1.760 ;
        RECT  5.175 0.770 5.335 1.760 ;
        RECT  4.045 0.770 5.175 0.930 ;
        RECT  4.875 0.380 5.135 0.590 ;
        RECT  4.835 1.140 4.995 2.100 ;
        RECT  3.705 0.430 4.875 0.590 ;
        RECT  4.545 1.140 4.835 1.300 ;
        RECT  4.495 1.620 4.655 2.560 ;
        RECT  4.225 1.620 4.495 1.780 ;
        RECT  3.025 2.400 4.495 2.560 ;
        RECT  4.045 1.990 4.285 2.150 ;
        RECT  3.885 0.770 4.045 2.150 ;
        RECT  3.395 0.990 3.885 1.190 ;
        RECT  3.545 0.430 3.705 0.810 ;
        RECT  3.095 0.650 3.545 0.810 ;
        RECT  3.095 1.495 3.495 1.755 ;
        RECT  2.755 0.310 3.365 0.470 ;
        RECT  2.935 0.650 3.095 2.175 ;
        RECT  2.865 2.355 3.025 2.560 ;
        RECT  1.445 2.015 2.935 2.175 ;
        RECT  1.105 2.355 2.865 2.515 ;
        RECT  2.595 0.310 2.755 1.835 ;
        RECT  1.825 1.675 2.595 1.835 ;
        RECT  1.825 0.755 1.895 0.915 ;
        RECT  1.665 0.755 1.825 1.835 ;
        RECT  1.530 0.310 1.790 0.575 ;
        RECT  1.635 0.755 1.665 0.915 ;
        RECT  1.635 1.675 1.665 1.835 ;
        RECT  0.945 0.415 1.530 0.575 ;
        RECT  1.285 1.765 1.445 2.175 ;
        RECT  1.285 0.755 1.385 0.915 ;
        RECT  1.125 0.755 1.285 1.570 ;
        RECT  1.105 1.410 1.125 1.570 ;
        RECT  0.945 1.410 1.105 2.515 ;
        RECT  0.785 0.415 0.945 0.865 ;
        RECT  0.385 0.705 0.785 0.865 ;
        RECT  0.285 0.705 0.385 0.965 ;
        RECT  0.285 1.915 0.385 2.175 ;
        RECT  0.125 0.705 0.285 2.175 ;
    END
END DFFHQNX4MTH

MACRO DFFHQNX8MTH
    CLASS CORE ;
    FOREIGN DFFHQNX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.525 1.935 9.185 2.435 ;
        RECT  8.525 0.810 9.045 1.010 ;
        RECT  7.995 0.810 8.525 2.435 ;
        RECT  7.805 0.810 7.995 1.010 ;
        END
        AntennaDiffArea 1.164 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 1.220 2.360 1.725 ;
        RECT  1.965 1.220 2.065 1.495 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.210 0.765 1.740 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.585 -0.130 10.250 0.130 ;
        RECT  9.325 -0.130 9.585 0.250 ;
        RECT  7.525 -0.130 9.325 0.130 ;
        RECT  7.265 -0.130 7.525 0.250 ;
        RECT  5.915 -0.130 7.265 0.130 ;
        RECT  5.315 -0.130 5.915 0.250 ;
        RECT  4.565 -0.130 5.315 0.130 ;
        RECT  3.625 -0.130 4.565 0.250 ;
        RECT  2.415 -0.130 3.625 0.130 ;
        RECT  2.215 -0.130 2.415 0.700 ;
        RECT  0.655 -0.130 2.215 0.130 ;
        RECT  0.395 -0.130 0.655 0.250 ;
        RECT  0.000 -0.130 0.395 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.715 2.740 10.250 3.000 ;
        RECT  6.775 2.570 7.715 3.000 ;
        RECT  5.855 2.740 6.775 3.000 ;
        RECT  4.915 2.620 5.855 3.000 ;
        RECT  0.765 2.740 4.915 3.000 ;
        RECT  0.165 2.455 0.765 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.125 0.425 10.155 1.735 ;
        RECT  9.995 0.425 10.125 2.375 ;
        RECT  9.865 0.425 9.995 0.925 ;
        RECT  9.865 1.575 9.995 2.375 ;
        RECT  9.315 1.575 9.865 1.735 ;
        RECT  9.675 1.135 9.785 1.395 ;
        RECT  9.515 0.430 9.675 1.395 ;
        RECT  7.535 0.430 9.515 0.590 ;
        RECT  9.155 1.260 9.315 1.735 ;
        RECT  8.705 1.260 9.155 1.520 ;
        RECT  7.375 0.430 7.535 2.070 ;
        RECT  6.995 0.430 7.375 0.590 ;
        RECT  6.855 1.910 7.375 2.070 ;
        RECT  6.915 1.445 7.175 1.705 ;
        RECT  6.735 0.355 6.995 0.590 ;
        RECT  6.555 1.445 6.915 1.605 ;
        RECT  6.595 1.910 6.855 2.170 ;
        RECT  6.415 0.430 6.555 1.605 ;
        RECT  6.425 2.400 6.515 2.560 ;
        RECT  6.165 2.280 6.425 2.560 ;
        RECT  6.395 0.350 6.415 1.605 ;
        RECT  6.155 0.350 6.395 0.590 ;
        RECT  5.745 0.990 6.215 1.150 ;
        RECT  5.745 1.940 6.210 2.100 ;
        RECT  4.625 2.280 6.165 2.440 ;
        RECT  4.980 0.430 6.155 0.590 ;
        RECT  5.585 0.990 5.745 2.100 ;
        RECT  4.965 1.940 5.585 2.100 ;
        RECT  5.305 1.600 5.405 1.760 ;
        RECT  5.145 0.770 5.305 1.760 ;
        RECT  4.045 0.770 5.145 0.930 ;
        RECT  4.720 0.380 4.980 0.590 ;
        RECT  4.805 1.140 4.965 2.100 ;
        RECT  4.535 1.140 4.805 1.300 ;
        RECT  3.705 0.430 4.720 0.590 ;
        RECT  4.465 1.620 4.625 2.560 ;
        RECT  4.225 1.620 4.465 1.780 ;
        RECT  3.025 2.400 4.465 2.560 ;
        RECT  4.045 1.990 4.285 2.150 ;
        RECT  3.885 0.770 4.045 2.150 ;
        RECT  3.395 0.990 3.885 1.190 ;
        RECT  3.545 0.430 3.705 0.810 ;
        RECT  3.095 0.650 3.545 0.810 ;
        RECT  3.095 1.495 3.495 1.755 ;
        RECT  2.755 0.310 3.365 0.470 ;
        RECT  2.935 0.650 3.095 2.175 ;
        RECT  2.865 2.355 3.025 2.560 ;
        RECT  1.445 2.015 2.935 2.175 ;
        RECT  1.105 2.355 2.865 2.515 ;
        RECT  2.595 0.310 2.755 1.040 ;
        RECT  1.895 0.880 2.595 1.040 ;
        RECT  1.785 0.755 1.895 1.040 ;
        RECT  1.785 1.675 1.885 1.835 ;
        RECT  1.530 0.310 1.790 0.575 ;
        RECT  1.625 0.755 1.785 1.835 ;
        RECT  0.945 0.415 1.530 0.575 ;
        RECT  1.285 1.765 1.445 2.175 ;
        RECT  1.285 0.755 1.385 0.915 ;
        RECT  1.125 0.755 1.285 1.410 ;
        RECT  1.105 1.250 1.125 1.410 ;
        RECT  0.945 1.250 1.105 2.515 ;
        RECT  0.785 0.415 0.945 0.865 ;
        RECT  0.385 0.705 0.785 0.865 ;
        RECT  0.285 0.705 0.385 0.965 ;
        RECT  0.285 1.915 0.385 2.175 ;
        RECT  0.125 0.705 0.285 2.175 ;
    END
END DFFHQNX8MTH

MACRO DFFHQX1MTH
    CLASS CORE ;
    FOREIGN DFFHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.690 8.920 1.990 ;
        RECT  8.635 0.690 8.710 0.950 ;
        RECT  8.635 1.730 8.710 1.990 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.440 1.370 ;
        RECT  2.085 1.105 2.150 1.370 ;
        END
        AntennaGateArea 0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.210 0.810 1.785 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.515 -0.130 9.020 0.130 ;
        RECT  7.575 -0.130 8.515 0.250 ;
        RECT  5.885 -0.130 7.575 0.130 ;
        RECT  5.285 -0.130 5.885 0.250 ;
        RECT  4.535 -0.130 5.285 0.130 ;
        RECT  4.275 -0.130 4.535 0.250 ;
        RECT  2.575 -0.130 4.275 0.130 ;
        RECT  2.315 -0.130 2.575 0.700 ;
        RECT  0.680 -0.130 2.315 0.130 ;
        RECT  0.520 -0.130 0.680 0.300 ;
        RECT  0.000 -0.130 0.520 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.515 2.740 9.020 3.000 ;
        RECT  7.575 2.570 8.515 3.000 ;
        RECT  5.725 2.740 7.575 3.000 ;
        RECT  4.785 2.620 5.725 3.000 ;
        RECT  4.465 2.740 4.785 3.000 ;
        RECT  3.525 2.620 4.465 3.000 ;
        RECT  3.210 2.740 3.525 3.000 ;
        RECT  2.270 2.620 3.210 3.000 ;
        RECT  0.860 2.740 2.270 3.000 ;
        RECT  0.260 2.620 0.860 3.000 ;
        RECT  0.000 2.740 0.260 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.265 1.260 8.365 1.520 ;
        RECT  8.105 0.430 8.265 2.310 ;
        RECT  6.895 0.430 8.105 0.590 ;
        RECT  6.895 2.150 8.105 2.310 ;
        RECT  7.665 0.770 7.925 1.965 ;
        RECT  7.575 0.770 7.665 0.930 ;
        RECT  7.515 1.235 7.665 1.495 ;
        RECT  7.135 1.500 7.235 1.660 ;
        RECT  6.975 1.145 7.135 1.660 ;
        RECT  6.555 1.145 6.975 1.305 ;
        RECT  6.735 0.365 6.895 0.965 ;
        RECT  6.735 1.870 6.895 2.470 ;
        RECT  6.555 1.495 6.690 1.655 ;
        RECT  6.445 0.430 6.555 1.305 ;
        RECT  6.395 1.495 6.555 2.440 ;
        RECT  6.395 0.335 6.445 1.305 ;
        RECT  6.185 0.335 6.395 0.590 ;
        RECT  4.920 2.280 6.395 2.440 ;
        RECT  6.055 0.770 6.215 2.090 ;
        RECT  3.215 0.430 6.185 0.590 ;
        RECT  5.310 1.655 6.055 1.815 ;
        RECT  5.775 1.215 5.875 1.475 ;
        RECT  5.615 0.820 5.775 1.475 ;
        RECT  4.360 0.820 5.615 0.980 ;
        RECT  5.150 1.430 5.310 1.815 ;
        RECT  4.760 1.485 4.920 2.440 ;
        RECT  4.730 1.485 4.760 1.645 ;
        RECT  1.150 2.280 4.760 2.440 ;
        RECT  4.570 1.385 4.730 1.645 ;
        RECT  4.360 1.825 4.580 2.085 ;
        RECT  4.200 0.770 4.360 2.085 ;
        RECT  3.395 0.770 4.200 0.930 ;
        RECT  3.720 1.110 3.880 2.100 ;
        RECT  3.215 1.110 3.720 1.270 ;
        RECT  1.490 1.940 3.720 2.100 ;
        RECT  3.190 1.450 3.450 1.760 ;
        RECT  3.055 0.430 3.215 1.270 ;
        RECT  1.905 1.600 3.190 1.760 ;
        RECT  2.885 0.630 3.055 0.890 ;
        RECT  1.905 0.680 1.970 0.840 ;
        RECT  1.745 0.680 1.905 1.760 ;
        RECT  1.600 0.310 1.860 0.500 ;
        RECT  1.710 0.680 1.745 0.840 ;
        RECT  1.020 0.340 1.600 0.500 ;
        RECT  1.330 1.545 1.490 2.100 ;
        RECT  1.360 0.680 1.460 0.840 ;
        RECT  1.200 0.680 1.360 1.340 ;
        RECT  1.150 1.180 1.200 1.340 ;
        RECT  0.990 1.180 1.150 2.440 ;
        RECT  0.860 0.340 1.020 0.790 ;
        RECT  0.405 0.630 0.860 0.790 ;
        RECT  0.330 0.630 0.405 0.890 ;
        RECT  0.330 1.965 0.385 2.125 ;
        RECT  0.170 0.630 0.330 2.125 ;
        RECT  0.125 1.965 0.170 2.125 ;
    END
END DFFHQX1MTH

MACRO DFFHQX2MTH
    CLASS CORE ;
    FOREIGN DFFHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.385 8.920 2.385 ;
        RECT  8.635 0.385 8.710 0.985 ;
        RECT  8.635 1.785 8.710 2.385 ;
        END
        AntennaDiffArea 0.521 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 0.880 2.360 1.420 ;
        RECT  2.005 1.110 2.105 1.420 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.145 0.765 1.715 ;
        END
        AntennaGateArea 0.1417 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 -0.130 9.020 0.130 ;
        RECT  7.360 -0.130 8.300 0.250 ;
        RECT  5.675 -0.130 7.360 0.130 ;
        RECT  5.415 -0.130 5.675 0.250 ;
        RECT  4.480 -0.130 5.415 0.130 ;
        RECT  4.220 -0.130 4.480 0.250 ;
        RECT  2.705 -0.130 4.220 0.130 ;
        RECT  2.445 -0.130 2.705 0.320 ;
        RECT  0.635 -0.130 2.445 0.130 ;
        RECT  0.475 -0.130 0.635 0.345 ;
        RECT  0.000 -0.130 0.475 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.320 2.740 9.020 3.000 ;
        RECT  7.720 2.570 8.320 3.000 ;
        RECT  6.080 2.740 7.720 3.000 ;
        RECT  5.820 2.620 6.080 3.000 ;
        RECT  4.995 2.740 5.820 3.000 ;
        RECT  4.735 2.620 4.995 3.000 ;
        RECT  3.400 2.740 4.735 3.000 ;
        RECT  3.140 2.620 3.400 3.000 ;
        RECT  2.445 2.740 3.140 3.000 ;
        RECT  2.185 2.620 2.445 3.000 ;
        RECT  0.765 2.740 2.185 3.000 ;
        RECT  0.225 2.425 0.765 3.000 ;
        RECT  0.000 2.740 0.225 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.330 1.205 8.400 1.465 ;
        RECT  8.170 0.430 8.330 2.235 ;
        RECT  6.995 0.430 8.170 0.590 ;
        RECT  7.075 2.075 8.170 2.235 ;
        RECT  7.695 0.770 7.955 1.895 ;
        RECT  7.665 0.770 7.695 1.495 ;
        RECT  7.555 1.235 7.665 1.495 ;
        RECT  6.555 1.475 7.275 1.635 ;
        RECT  6.815 1.855 7.075 2.455 ;
        RECT  6.735 0.355 6.995 0.590 ;
        RECT  5.895 1.845 6.565 2.005 ;
        RECT  6.395 0.430 6.555 1.635 ;
        RECT  5.070 0.430 6.395 0.590 ;
        RECT  6.155 1.155 6.395 1.365 ;
        RECT  6.045 2.215 6.305 2.440 ;
        RECT  5.895 0.785 6.215 0.945 ;
        RECT  4.595 2.280 6.045 2.440 ;
        RECT  5.735 0.785 5.895 2.100 ;
        RECT  4.935 1.940 5.735 2.100 ;
        RECT  5.495 1.570 5.545 1.730 ;
        RECT  5.335 0.770 5.495 1.730 ;
        RECT  3.895 0.770 5.335 0.930 ;
        RECT  5.285 1.570 5.335 1.730 ;
        RECT  4.810 0.335 5.070 0.590 ;
        RECT  4.775 1.255 4.935 2.100 ;
        RECT  4.040 0.430 4.810 0.590 ;
        RECT  4.675 1.255 4.775 1.415 ;
        RECT  4.435 1.600 4.595 2.440 ;
        RECT  4.395 1.600 4.435 1.760 ;
        RECT  1.105 2.280 4.435 2.440 ;
        RECT  4.135 1.570 4.395 1.760 ;
        RECT  3.895 1.940 4.255 2.100 ;
        RECT  3.880 0.310 4.040 0.590 ;
        RECT  3.735 0.770 3.895 2.100 ;
        RECT  3.105 0.310 3.880 0.470 ;
        RECT  3.600 0.770 3.735 0.930 ;
        RECT  3.340 0.650 3.600 0.930 ;
        RECT  3.395 1.110 3.555 2.100 ;
        RECT  3.105 1.110 3.395 1.270 ;
        RECT  1.445 1.940 3.395 2.100 ;
        RECT  3.025 1.540 3.125 1.700 ;
        RECT  2.945 0.310 3.105 1.270 ;
        RECT  2.865 1.540 3.025 1.760 ;
        RECT  2.880 0.570 2.945 0.830 ;
        RECT  1.785 1.600 2.865 1.760 ;
        RECT  2.700 1.010 2.765 1.270 ;
        RECT  2.540 0.540 2.700 1.270 ;
        RECT  2.265 0.540 2.540 0.700 ;
        RECT  2.105 0.310 2.265 0.700 ;
        RECT  0.975 0.310 2.105 0.470 ;
        RECT  1.785 0.680 1.925 0.840 ;
        RECT  1.625 0.680 1.785 1.760 ;
        RECT  1.285 1.665 1.445 2.100 ;
        RECT  1.365 0.680 1.415 0.840 ;
        RECT  1.205 0.680 1.365 1.230 ;
        RECT  1.155 0.680 1.205 0.840 ;
        RECT  1.105 1.070 1.205 1.230 ;
        RECT  0.945 1.070 1.105 2.440 ;
        RECT  0.815 0.310 0.975 0.865 ;
        RECT  0.335 0.705 0.815 0.865 ;
        RECT  0.285 1.895 0.385 2.055 ;
        RECT  0.285 0.705 0.335 0.965 ;
        RECT  0.125 0.705 0.285 2.055 ;
    END
END DFFHQX2MTH

MACRO DFFHQX4MTH
    CLASS CORE ;
    FOREIGN DFFHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.705 1.290 9.740 1.580 ;
        RECT  9.445 0.400 9.705 2.380 ;
        END
        AntennaDiffArea 0.582 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.280 2.030 1.490 ;
        RECT  1.330 1.280 1.540 1.580 ;
        END
        AntennaGateArea 0.0806 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.650 1.190 0.810 1.785 ;
        RECT  0.465 1.190 0.650 1.580 ;
        END
        AntennaGateArea 0.2158 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.195 -0.130 10.250 0.130 ;
        RECT  8.935 -0.130 9.195 1.025 ;
        RECT  8.905 -0.130 8.935 0.250 ;
        RECT  8.385 -0.130 8.905 0.130 ;
        RECT  7.785 -0.130 8.385 0.250 ;
        RECT  6.105 -0.130 7.785 0.130 ;
        RECT  5.505 -0.130 6.105 0.250 ;
        RECT  4.805 -0.130 5.505 0.130 ;
        RECT  4.545 -0.130 4.805 0.250 ;
        RECT  2.405 -0.130 4.545 0.130 ;
        RECT  2.145 -0.130 2.405 0.755 ;
        RECT  0.510 -0.130 2.145 0.130 ;
        RECT  0.250 -0.130 0.510 0.250 ;
        RECT  0.000 -0.130 0.250 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.165 2.740 10.250 3.000 ;
        RECT  8.565 2.415 9.165 3.000 ;
        RECT  5.195 2.740 8.565 3.000 ;
        RECT  4.595 2.570 5.195 3.000 ;
        RECT  3.505 2.740 4.595 3.000 ;
        RECT  3.345 2.570 3.505 3.000 ;
        RECT  0.785 2.740 3.345 3.000 ;
        RECT  0.185 2.260 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.100 1.210 9.200 1.470 ;
        RECT  8.940 1.210 9.100 2.235 ;
        RECT  7.785 2.075 8.940 2.235 ;
        RECT  8.525 1.735 8.735 1.895 ;
        RECT  8.525 0.765 8.625 1.025 ;
        RECT  8.265 0.765 8.525 1.895 ;
        RECT  7.945 1.530 8.045 1.690 ;
        RECT  7.785 0.430 7.945 1.690 ;
        RECT  7.525 0.430 7.785 0.590 ;
        RECT  7.695 1.945 7.785 2.445 ;
        RECT  7.585 1.945 7.695 2.560 ;
        RECT  7.405 0.770 7.585 2.560 ;
        RECT  7.265 0.310 7.525 0.590 ;
        RECT  6.895 0.770 7.405 0.930 ;
        RECT  6.765 2.400 7.405 2.560 ;
        RECT  4.170 0.430 7.265 0.590 ;
        RECT  7.135 1.880 7.225 2.140 ;
        RECT  6.975 1.110 7.135 2.140 ;
        RECT  6.645 1.110 6.975 1.270 ;
        RECT  6.555 2.285 6.765 2.560 ;
        RECT  6.385 0.820 6.645 1.270 ;
        RECT  6.505 2.285 6.555 2.445 ;
        RECT  6.295 1.475 6.455 2.110 ;
        RECT  6.035 1.110 6.385 1.270 ;
        RECT  6.100 1.950 6.295 2.110 ;
        RECT  5.940 1.950 6.100 2.390 ;
        RECT  5.875 1.110 6.035 1.765 ;
        RECT  4.695 2.230 5.940 2.390 ;
        RECT  5.735 1.605 5.875 1.765 ;
        RECT  5.475 1.605 5.735 2.050 ;
        RECT  5.505 0.815 5.665 1.425 ;
        RECT  4.055 0.815 5.505 0.975 ;
        RECT  5.035 1.605 5.475 1.765 ;
        RECT  4.875 1.365 5.035 1.765 ;
        RECT  4.535 1.245 4.695 2.390 ;
        RECT  4.345 1.245 4.535 1.505 ;
        RECT  4.425 2.130 4.535 2.390 ;
        RECT  3.055 2.130 4.425 2.290 ;
        RECT  4.055 1.685 4.355 1.945 ;
        RECT  4.010 0.390 4.170 0.590 ;
        RECT  3.955 0.815 4.055 1.945 ;
        RECT  3.515 0.390 4.010 0.550 ;
        RECT  3.895 0.765 3.955 1.945 ;
        RECT  3.695 0.765 3.895 1.025 ;
        RECT  3.105 1.290 3.705 1.550 ;
        RECT  3.355 0.390 3.515 0.875 ;
        RECT  3.100 0.715 3.355 0.875 ;
        RECT  2.760 0.310 3.175 0.470 ;
        RECT  3.100 1.290 3.105 1.895 ;
        RECT  2.940 0.715 3.100 1.895 ;
        RECT  2.895 2.130 3.055 2.560 ;
        RECT  2.710 1.735 2.940 1.895 ;
        RECT  1.585 2.400 2.895 2.560 ;
        RECT  2.600 0.310 2.760 1.095 ;
        RECT  2.550 1.735 2.710 2.220 ;
        RECT  2.370 0.935 2.600 1.095 ;
        RECT  1.765 2.060 2.550 2.220 ;
        RECT  2.210 0.935 2.370 1.850 ;
        RECT  1.835 0.935 2.210 1.095 ;
        RECT  1.905 1.690 2.210 1.850 ;
        RECT  1.675 0.715 1.835 1.095 ;
        RECT  0.850 0.310 1.725 0.470 ;
        RECT  1.575 0.715 1.675 0.875 ;
        RECT  1.150 1.760 1.585 2.560 ;
        RECT  1.150 0.730 1.325 0.890 ;
        RECT  0.990 0.730 1.150 2.560 ;
        RECT  0.690 0.310 0.850 0.590 ;
        RECT  0.385 0.430 0.690 0.590 ;
        RECT  0.285 0.430 0.385 1.010 ;
        RECT  0.285 1.760 0.385 1.920 ;
        RECT  0.125 0.430 0.285 1.920 ;
    END
END DFFHQX4MTH

MACRO DFFHQX8MTH
    CLASS CORE ;
    FOREIGN DFFHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.965 0.400 11.225 2.380 ;
        RECT  10.145 1.075 10.965 1.795 ;
        RECT  9.895 0.400 10.145 2.380 ;
        END
        AntennaDiffArea 1.164 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.280 2.440 1.540 ;
        RECT  1.880 1.280 2.110 1.455 ;
        END
        AntennaGateArea 0.1534 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.175 0.800 1.625 ;
        END
        AntennaGateArea 0.2925 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 -0.130 11.890 0.130 ;
        RECT  11.505 -0.130 11.765 0.980 ;
        RECT  10.685 -0.130 11.505 0.130 ;
        RECT  10.425 -0.130 10.685 0.805 ;
        RECT  9.625 -0.130 10.425 0.130 ;
        RECT  9.365 -0.130 9.625 0.975 ;
        RECT  8.795 -0.130 9.365 0.130 ;
        RECT  8.195 -0.130 8.795 0.250 ;
        RECT  6.515 -0.130 8.195 0.130 ;
        RECT  5.915 -0.130 6.515 0.250 ;
        RECT  5.045 -0.130 5.915 0.130 ;
        RECT  4.785 -0.130 5.045 0.250 ;
        RECT  2.515 -0.130 4.785 0.130 ;
        RECT  2.255 -0.130 2.515 0.250 ;
        RECT  1.265 -0.130 2.255 0.130 ;
        RECT  0.665 -0.130 1.265 0.250 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 2.740 11.890 3.000 ;
        RECT  11.505 1.890 11.765 3.000 ;
        RECT  10.685 2.740 11.505 3.000 ;
        RECT  10.425 2.015 10.685 3.000 ;
        RECT  9.425 2.740 10.425 3.000 ;
        RECT  8.825 2.465 9.425 3.000 ;
        RECT  6.575 2.740 8.825 3.000 ;
        RECT  6.315 2.570 6.575 3.000 ;
        RECT  5.495 2.740 6.315 3.000 ;
        RECT  4.895 2.570 5.495 3.000 ;
        RECT  3.805 2.740 4.895 3.000 ;
        RECT  3.645 2.570 3.805 3.000 ;
        RECT  0.795 2.740 3.645 3.000 ;
        RECT  0.195 2.475 0.795 3.000 ;
        RECT  0.000 2.740 0.195 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.345 1.205 9.715 1.465 ;
        RECT  9.185 1.205 9.345 2.285 ;
        RECT  8.105 2.125 9.185 2.285 ;
        RECT  8.945 0.765 9.055 1.025 ;
        RECT  8.945 1.685 9.005 1.945 ;
        RECT  8.685 0.765 8.945 1.945 ;
        RECT  8.585 1.315 8.685 1.575 ;
        RECT  8.205 0.430 8.365 1.735 ;
        RECT  7.935 0.430 8.205 0.590 ;
        RECT  8.105 1.575 8.205 1.735 ;
        RECT  7.885 1.945 8.105 2.560 ;
        RECT  7.675 0.310 7.935 0.590 ;
        RECT  7.725 0.770 7.885 2.560 ;
        RECT  7.305 0.770 7.725 0.930 ;
        RECT  7.095 2.400 7.725 2.560 ;
        RECT  4.580 0.430 7.675 0.590 ;
        RECT  7.385 1.110 7.545 2.140 ;
        RECT  7.055 1.110 7.385 1.270 ;
        RECT  6.875 2.235 7.095 2.560 ;
        RECT  6.795 0.770 7.055 1.270 ;
        RECT  6.385 1.110 6.795 1.270 ;
        RECT  6.730 1.500 6.775 1.760 ;
        RECT  6.570 1.500 6.730 2.110 ;
        RECT  6.400 1.950 6.570 2.110 ;
        RECT  6.240 1.950 6.400 2.390 ;
        RECT  6.225 1.110 6.385 1.765 ;
        RECT  4.995 2.230 6.240 2.390 ;
        RECT  6.035 1.605 6.225 1.765 ;
        RECT  5.785 0.815 6.045 1.425 ;
        RECT  5.775 1.605 6.035 2.050 ;
        RECT  4.375 0.815 5.785 0.975 ;
        RECT  5.335 1.605 5.775 1.765 ;
        RECT  5.175 1.365 5.335 1.765 ;
        RECT  4.835 1.245 4.995 2.390 ;
        RECT  4.645 1.245 4.835 1.505 ;
        RECT  3.465 2.140 4.835 2.300 ;
        RECT  4.375 1.695 4.655 1.955 ;
        RECT  4.420 0.380 4.580 0.590 ;
        RECT  3.805 0.380 4.420 0.540 ;
        RECT  4.215 0.815 4.375 1.955 ;
        RECT  4.145 0.815 4.215 1.025 ;
        RECT  3.985 0.765 4.145 1.025 ;
        RECT  3.635 1.290 4.035 1.550 ;
        RECT  3.645 0.380 3.805 0.910 ;
        RECT  3.635 0.750 3.645 0.910 ;
        RECT  3.475 0.750 3.635 1.905 ;
        RECT  3.120 1.745 3.475 1.905 ;
        RECT  3.295 0.310 3.465 0.570 ;
        RECT  3.305 2.140 3.465 2.560 ;
        RECT  1.595 2.400 3.305 2.560 ;
        RECT  3.135 0.310 3.295 1.095 ;
        RECT  2.780 0.935 3.135 1.095 ;
        RECT  2.960 1.745 3.120 2.220 ;
        RECT  1.935 2.060 2.960 2.220 ;
        RECT  2.695 0.310 2.955 0.590 ;
        RECT  2.620 0.935 2.780 1.880 ;
        RECT  0.385 0.430 2.695 0.590 ;
        RECT  1.975 0.935 2.620 1.095 ;
        RECT  2.115 1.720 2.620 1.880 ;
        RECT  1.715 0.800 1.975 1.095 ;
        RECT  1.775 1.635 1.935 2.220 ;
        RECT  1.600 1.635 1.775 1.795 ;
        RECT  1.340 1.455 1.600 1.795 ;
        RECT  1.435 1.975 1.595 2.560 ;
        RECT  1.140 0.800 1.455 0.960 ;
        RECT  1.140 1.975 1.435 2.135 ;
        RECT  0.980 0.800 1.140 2.135 ;
        RECT  0.285 0.430 0.385 1.010 ;
        RECT  0.285 1.825 0.385 2.085 ;
        RECT  0.125 0.430 0.285 2.085 ;
    END
END DFFHQX8MTH

MACRO DFFHX1MTH
    CLASS CORE ;
    FOREIGN DFFHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.940 0.765 10.150 1.995 ;
        RECT  9.865 0.765 9.940 1.025 ;
        RECT  9.835 1.735 9.940 1.995 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.815 8.920 1.995 ;
        END
        AntennaDiffArea 0.289 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.145 2.435 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.145 0.355 1.895 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.925 -0.130 10.250 0.130 ;
        RECT  9.645 -0.130 9.925 0.300 ;
        RECT  9.450 -0.130 9.645 0.130 ;
        RECT  8.950 -0.130 9.450 0.300 ;
        RECT  8.030 -0.130 8.950 0.130 ;
        RECT  7.870 -0.130 8.030 0.620 ;
        RECT  6.280 -0.130 7.870 0.130 ;
        RECT  6.020 -0.130 6.280 0.250 ;
        RECT  5.120 -0.130 6.020 0.130 ;
        RECT  4.860 -0.130 5.120 0.250 ;
        RECT  0.355 -0.130 4.860 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.800 2.740 10.250 3.000 ;
        RECT  9.300 2.570 9.800 3.000 ;
        RECT  8.190 2.740 9.300 3.000 ;
        RECT  8.030 2.245 8.190 3.000 ;
        RECT  5.770 2.740 8.030 3.000 ;
        RECT  5.170 2.205 5.770 3.000 ;
        RECT  4.365 2.740 5.170 3.000 ;
        RECT  3.425 2.620 4.365 3.000 ;
        RECT  2.975 2.740 3.425 3.000 ;
        RECT  2.035 2.620 2.975 3.000 ;
        RECT  0.810 2.740 2.035 3.000 ;
        RECT  0.550 2.620 0.810 3.000 ;
        RECT  0.000 2.740 0.550 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.260 1.250 9.705 1.510 ;
        RECT  9.100 1.250 9.260 2.335 ;
        RECT  8.940 2.175 9.100 2.335 ;
        RECT  8.680 2.175 8.940 2.560 ;
        RECT  8.530 2.175 8.680 2.335 ;
        RECT  8.530 0.355 8.650 0.565 ;
        RECT  8.370 0.355 8.530 2.335 ;
        RECT  8.000 1.265 8.370 1.525 ;
        RECT  7.480 2.400 7.850 2.560 ;
        RECT  7.670 0.810 7.730 1.710 ;
        RECT  7.570 0.435 7.670 1.710 ;
        RECT  7.510 0.435 7.570 0.975 ;
        RECT  7.160 0.435 7.510 0.595 ;
        RECT  7.380 1.955 7.480 2.560 ;
        RECT  7.330 1.185 7.380 2.560 ;
        RECT  7.220 0.815 7.330 2.560 ;
        RECT  7.170 0.815 7.220 1.345 ;
        RECT  7.070 0.815 7.170 0.975 ;
        RECT  6.900 0.345 7.160 0.595 ;
        RECT  6.850 1.840 6.920 2.100 ;
        RECT  5.680 0.435 6.900 0.595 ;
        RECT  6.690 0.800 6.850 2.100 ;
        RECT  6.240 2.385 6.710 2.545 ;
        RECT  6.560 0.800 6.690 0.960 ;
        RECT  6.420 1.525 6.690 2.100 ;
        RECT  6.310 1.185 6.480 1.345 ;
        RECT  5.220 1.525 6.420 1.685 ;
        RECT  6.150 0.800 6.310 1.345 ;
        RECT  6.080 1.865 6.240 2.545 ;
        RECT  4.210 0.800 6.150 0.960 ;
        RECT  4.910 1.865 6.080 2.025 ;
        RECT  5.420 0.325 5.680 0.595 ;
        RECT  4.555 0.435 5.420 0.595 ;
        RECT  5.060 1.195 5.220 1.685 ;
        RECT  4.960 1.195 5.060 1.355 ;
        RECT  4.860 1.865 4.910 2.505 ;
        RECT  4.750 1.865 4.860 2.560 ;
        RECT  4.700 2.250 4.750 2.560 ;
        RECT  1.695 2.250 4.700 2.410 ;
        RECT  4.395 0.380 4.555 0.595 ;
        RECT  4.210 1.690 4.485 1.950 ;
        RECT  3.870 0.380 4.395 0.540 ;
        RECT  4.050 0.720 4.210 1.950 ;
        RECT  3.710 0.380 3.870 0.910 ;
        RECT  3.685 1.290 3.835 1.550 ;
        RECT  3.685 0.750 3.710 0.910 ;
        RECT  3.525 0.750 3.685 2.070 ;
        RECT  3.370 0.310 3.530 0.570 ;
        RECT  3.455 0.750 3.525 1.010 ;
        RECT  1.445 1.910 3.525 2.070 ;
        RECT  3.275 0.410 3.370 0.570 ;
        RECT  3.115 0.410 3.275 0.810 ;
        RECT  1.925 0.650 3.115 0.810 ;
        RECT  0.695 0.310 2.935 0.470 ;
        RECT  1.765 0.650 1.925 1.730 ;
        RECT  1.675 0.650 1.765 0.810 ;
        RECT  1.665 1.570 1.765 1.730 ;
        RECT  1.435 2.250 1.695 2.510 ;
        RECT  1.445 1.020 1.495 1.180 ;
        RECT  1.285 0.990 1.445 2.070 ;
        RECT  1.035 2.250 1.435 2.410 ;
        RECT  1.035 0.650 1.425 0.810 ;
        RECT  1.235 1.020 1.285 1.180 ;
        RECT  0.875 0.650 1.035 2.410 ;
        RECT  0.535 0.310 0.695 2.250 ;
        RECT  0.125 0.700 0.535 0.960 ;
        RECT  0.385 2.090 0.535 2.250 ;
        RECT  0.125 2.090 0.385 2.350 ;
    END
END DFFHX1MTH

MACRO DFFHX2MTH
    CLASS CORE ;
    FOREIGN DFFHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.305 0.765 10.560 1.950 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.290 1.290 9.330 1.580 ;
        RECT  9.180 0.425 9.290 1.580 ;
        RECT  9.020 0.425 9.180 1.985 ;
        END
        AntennaDiffArea 0.417 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.470 1.755 1.950 ;
        END
        AntennaGateArea 0.0923 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.355 1.910 ;
        END
        AntennaGateArea 0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.170 -0.130 10.660 0.130 ;
        RECT  9.830 -0.130 10.170 0.300 ;
        RECT  9.570 -0.130 9.830 1.025 ;
        RECT  8.080 -0.130 9.570 0.130 ;
        RECT  7.820 -0.130 8.080 0.250 ;
        RECT  6.280 -0.130 7.820 0.130 ;
        RECT  6.020 -0.130 6.280 0.250 ;
        RECT  5.120 -0.130 6.020 0.130 ;
        RECT  4.860 -0.130 5.120 0.250 ;
        RECT  2.635 -0.130 4.860 0.130 ;
        RECT  2.375 -0.130 2.635 0.250 ;
        RECT  0.355 -0.130 2.375 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.110 2.740 10.660 3.000 ;
        RECT  9.850 2.170 10.110 3.000 ;
        RECT  9.510 2.570 9.850 3.000 ;
        RECT  8.480 2.740 9.510 3.000 ;
        RECT  8.320 2.235 8.480 3.000 ;
        RECT  5.280 2.740 8.320 3.000 ;
        RECT  5.020 2.620 5.280 3.000 ;
        RECT  0.810 2.740 5.020 3.000 ;
        RECT  0.210 2.570 0.810 3.000 ;
        RECT  0.000 2.740 0.210 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.835 1.250 10.095 1.510 ;
        RECT  9.670 1.350 9.835 1.510 ;
        RECT  9.510 1.350 9.670 2.325 ;
        RECT  9.260 2.165 9.510 2.325 ;
        RECT  9.000 2.165 9.260 2.515 ;
        RECT  8.820 2.165 9.000 2.325 ;
        RECT  8.660 1.265 8.820 2.325 ;
        RECT  8.650 1.265 8.660 1.525 ;
        RECT  8.390 0.440 8.650 1.525 ;
        RECT  8.320 1.265 8.390 1.525 ;
        RECT  7.840 2.400 8.140 2.560 ;
        RECT  7.890 0.435 8.050 1.715 ;
        RECT  7.590 0.435 7.890 0.595 ;
        RECT  7.630 1.940 7.840 2.560 ;
        RECT  7.620 1.940 7.630 2.100 ;
        RECT  6.940 2.400 7.630 2.560 ;
        RECT  7.460 0.815 7.620 2.100 ;
        RECT  7.330 0.310 7.590 0.595 ;
        RECT  7.070 0.815 7.460 0.975 ;
        RECT  5.680 0.435 7.330 0.595 ;
        RECT  7.120 1.525 7.280 2.075 ;
        RECT  6.850 1.525 7.120 1.690 ;
        RECT  6.780 1.875 6.940 2.560 ;
        RECT  6.690 0.800 6.850 1.690 ;
        RECT  6.480 1.875 6.780 2.035 ;
        RECT  6.560 0.800 6.690 0.960 ;
        RECT  5.830 1.530 6.690 1.690 ;
        RECT  6.340 2.230 6.600 2.545 ;
        RECT  6.310 1.190 6.480 1.350 ;
        RECT  4.840 2.230 6.340 2.390 ;
        RECT  6.150 0.820 6.310 1.350 ;
        RECT  4.210 0.820 6.150 0.980 ;
        RECT  5.570 1.530 5.830 2.050 ;
        RECT  5.420 0.325 5.680 0.595 ;
        RECT  5.220 1.530 5.570 1.690 ;
        RECT  4.555 0.435 5.420 0.595 ;
        RECT  5.060 1.195 5.220 1.690 ;
        RECT  4.960 1.195 5.060 1.355 ;
        RECT  4.580 2.230 4.840 2.560 ;
        RECT  1.665 2.400 4.580 2.560 ;
        RECT  4.395 0.380 4.555 0.595 ;
        RECT  3.870 0.380 4.395 0.540 ;
        RECT  4.210 1.690 4.385 1.950 ;
        RECT  4.050 0.720 4.210 1.950 ;
        RECT  3.735 0.380 3.870 1.010 ;
        RECT  3.710 0.380 3.735 1.550 ;
        RECT  3.635 0.750 3.710 1.550 ;
        RECT  3.540 0.750 3.635 2.120 ;
        RECT  3.475 1.290 3.540 2.120 ;
        RECT  3.345 0.310 3.530 0.570 ;
        RECT  3.085 1.960 3.475 2.120 ;
        RECT  3.185 0.310 3.345 1.110 ;
        RECT  2.475 0.950 3.185 1.110 ;
        RECT  2.825 1.960 3.085 2.220 ;
        RECT  2.845 0.350 3.005 0.610 ;
        RECT  2.195 0.450 2.845 0.610 ;
        RECT  2.095 2.060 2.825 2.220 ;
        RECT  2.475 1.670 2.575 1.880 ;
        RECT  2.315 0.790 2.475 1.880 ;
        RECT  1.845 0.790 2.315 0.950 ;
        RECT  2.035 0.310 2.195 0.610 ;
        RECT  1.935 1.130 2.095 2.220 ;
        RECT  0.695 0.310 2.035 0.470 ;
        RECT  1.495 1.130 1.935 1.290 ;
        RECT  1.685 0.650 1.845 0.950 ;
        RECT  1.405 2.130 1.665 2.560 ;
        RECT  1.235 1.040 1.495 1.290 ;
        RECT  1.035 2.130 1.405 2.290 ;
        RECT  1.035 0.670 1.385 0.830 ;
        RECT  0.875 0.670 1.035 2.290 ;
        RECT  0.535 0.310 0.695 2.250 ;
        RECT  0.125 0.765 0.535 1.025 ;
        RECT  0.385 2.090 0.535 2.250 ;
        RECT  0.125 2.090 0.385 2.325 ;
    END
END DFFHX2MTH

MACRO DFFHX4MTH
    CLASS CORE ;
    FOREIGN DFFHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.760 0.765 10.970 1.945 ;
        RECT  10.685 0.765 10.760 1.025 ;
        RECT  10.685 1.685 10.760 1.945 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.965 1.290 10.150 1.580 ;
        RECT  9.710 0.425 9.965 1.945 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.530 1.755 1.990 ;
        END
        AntennaGateArea 0.1586 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.210 0.355 1.840 ;
        END
        AntennaGateArea 0.2041 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.505 -0.130 11.070 0.130 ;
        RECT  10.245 -0.130 10.505 0.570 ;
        RECT  9.455 -0.130 10.245 0.130 ;
        RECT  9.195 -0.130 9.455 1.020 ;
        RECT  8.325 -0.130 9.195 0.130 ;
        RECT  8.165 -0.130 8.325 0.730 ;
        RECT  6.280 -0.130 8.165 0.130 ;
        RECT  6.020 -0.130 6.280 0.250 ;
        RECT  5.120 -0.130 6.020 0.130 ;
        RECT  4.860 -0.130 5.120 0.250 ;
        RECT  0.355 -0.130 4.860 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.505 2.740 11.070 3.000 ;
        RECT  10.245 2.465 10.505 3.000 ;
        RECT  9.425 2.740 10.245 3.000 ;
        RECT  9.165 2.465 9.425 3.000 ;
        RECT  8.805 2.740 9.165 3.000 ;
        RECT  8.545 2.465 8.805 3.000 ;
        RECT  5.280 2.740 8.545 3.000 ;
        RECT  5.020 2.620 5.280 3.000 ;
        RECT  0.830 2.740 5.020 3.000 ;
        RECT  0.555 2.620 0.830 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.500 1.245 10.580 1.505 ;
        RECT  10.340 1.245 10.500 2.285 ;
        RECT  9.515 2.125 10.340 2.285 ;
        RECT  9.355 1.785 9.515 2.285 ;
        RECT  8.975 1.785 9.355 1.945 ;
        RECT  7.865 2.125 9.175 2.285 ;
        RECT  8.945 1.685 8.975 1.945 ;
        RECT  8.715 0.490 8.945 1.945 ;
        RECT  8.685 0.490 8.715 1.400 ;
        RECT  8.345 1.135 8.685 1.400 ;
        RECT  7.985 1.450 8.075 1.710 ;
        RECT  7.825 0.435 7.985 1.710 ;
        RECT  7.645 1.900 7.865 2.500 ;
        RECT  7.615 0.435 7.825 0.595 ;
        RECT  7.485 0.815 7.645 2.500 ;
        RECT  7.355 0.310 7.615 0.595 ;
        RECT  7.070 0.815 7.485 0.975 ;
        RECT  6.965 2.340 7.485 2.500 ;
        RECT  5.680 0.435 7.355 0.595 ;
        RECT  7.145 1.525 7.305 2.075 ;
        RECT  6.850 1.525 7.145 1.715 ;
        RECT  6.805 1.895 6.965 2.500 ;
        RECT  6.690 0.800 6.850 1.715 ;
        RECT  6.505 1.895 6.805 2.055 ;
        RECT  6.560 0.800 6.690 0.960 ;
        RECT  5.830 1.555 6.690 1.715 ;
        RECT  6.365 2.235 6.625 2.550 ;
        RECT  6.310 1.215 6.480 1.375 ;
        RECT  4.840 2.235 6.365 2.395 ;
        RECT  6.150 0.820 6.310 1.375 ;
        RECT  4.465 0.820 6.150 0.980 ;
        RECT  5.570 1.555 5.830 2.050 ;
        RECT  5.420 0.325 5.680 0.595 ;
        RECT  5.220 1.555 5.570 1.715 ;
        RECT  4.555 0.435 5.420 0.595 ;
        RECT  5.060 1.195 5.220 1.715 ;
        RECT  4.960 1.195 5.060 1.355 ;
        RECT  4.580 2.235 4.840 2.560 ;
        RECT  1.665 2.400 4.580 2.560 ;
        RECT  4.395 0.380 4.555 0.595 ;
        RECT  4.305 0.820 4.465 1.950 ;
        RECT  3.870 0.380 4.395 0.540 ;
        RECT  4.210 0.820 4.305 0.980 ;
        RECT  4.050 0.720 4.210 0.980 ;
        RECT  3.815 0.380 3.870 0.910 ;
        RECT  3.710 0.380 3.815 2.220 ;
        RECT  3.655 0.750 3.710 2.220 ;
        RECT  3.455 0.750 3.655 1.010 ;
        RECT  2.095 2.060 3.655 2.220 ;
        RECT  3.275 0.310 3.530 0.470 ;
        RECT  3.115 0.310 3.275 0.810 ;
        RECT  2.635 0.650 3.115 0.810 ;
        RECT  0.695 0.310 2.935 0.470 ;
        RECT  2.475 0.650 2.635 1.880 ;
        RECT  1.625 0.650 2.475 0.810 ;
        RECT  2.375 1.720 2.475 1.880 ;
        RECT  1.935 1.110 2.095 2.220 ;
        RECT  1.485 1.110 1.935 1.270 ;
        RECT  1.405 2.170 1.665 2.560 ;
        RECT  1.150 2.170 1.405 2.330 ;
        RECT  1.150 0.735 1.305 0.995 ;
        RECT  0.990 0.735 1.150 2.330 ;
        RECT  0.535 0.310 0.695 2.180 ;
        RECT  0.125 0.750 0.535 1.010 ;
        RECT  0.385 2.020 0.535 2.180 ;
        RECT  0.125 2.020 0.385 2.280 ;
    END
END DFFHX4MTH

MACRO DFFHX8MTH
    CLASS CORE ;
    FOREIGN DFFHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.580 0.765 11.790 1.945 ;
        RECT  11.505 0.765 11.580 1.025 ;
        RECT  11.505 1.685 11.580 1.945 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.540 0.425 10.795 1.945 ;
        RECT  9.865 1.290 10.540 1.580 ;
        RECT  9.610 0.425 9.865 1.945 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.530 1.755 1.990 ;
        END
        AntennaGateArea 0.1586 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.210 0.355 1.840 ;
        END
        AntennaGateArea 0.2041 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.335 -0.130 11.890 0.130 ;
        RECT  11.075 -0.130 11.335 0.570 ;
        RECT  9.325 -0.130 11.075 0.130 ;
        RECT  9.065 -0.130 9.325 0.385 ;
        RECT  8.325 -0.130 9.065 0.130 ;
        RECT  8.165 -0.130 8.325 0.730 ;
        RECT  6.280 -0.130 8.165 0.130 ;
        RECT  6.020 -0.130 6.280 0.250 ;
        RECT  5.120 -0.130 6.020 0.130 ;
        RECT  4.860 -0.130 5.120 0.250 ;
        RECT  0.355 -0.130 4.860 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.335 2.740 11.890 3.000 ;
        RECT  11.075 2.465 11.335 3.000 ;
        RECT  9.255 2.740 11.075 3.000 ;
        RECT  8.655 2.530 9.255 3.000 ;
        RECT  5.280 2.740 8.655 3.000 ;
        RECT  5.020 2.620 5.280 3.000 ;
        RECT  0.830 2.740 5.020 3.000 ;
        RECT  0.555 2.620 0.830 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.320 1.245 11.400 1.505 ;
        RECT  11.160 1.245 11.320 2.285 ;
        RECT  9.415 2.125 11.160 2.285 ;
        RECT  9.255 1.785 9.415 2.285 ;
        RECT  8.945 1.785 9.255 1.945 ;
        RECT  7.840 2.125 9.075 2.285 ;
        RECT  8.685 0.685 8.945 1.945 ;
        RECT  8.615 1.310 8.685 1.945 ;
        RECT  8.345 1.310 8.615 1.575 ;
        RECT  7.960 1.625 8.075 1.885 ;
        RECT  7.800 0.435 7.960 1.885 ;
        RECT  7.620 2.125 7.840 2.385 ;
        RECT  7.590 0.435 7.800 0.595 ;
        RECT  7.460 0.815 7.620 2.385 ;
        RECT  7.330 0.310 7.590 0.595 ;
        RECT  7.070 0.815 7.460 0.975 ;
        RECT  6.940 2.225 7.460 2.385 ;
        RECT  5.680 0.435 7.330 0.595 ;
        RECT  7.120 1.525 7.280 2.045 ;
        RECT  6.850 1.525 7.120 1.715 ;
        RECT  6.780 1.895 6.940 2.385 ;
        RECT  6.690 0.800 6.850 1.715 ;
        RECT  6.480 1.895 6.780 2.055 ;
        RECT  6.560 0.800 6.690 0.960 ;
        RECT  5.830 1.555 6.690 1.715 ;
        RECT  6.340 2.235 6.600 2.550 ;
        RECT  6.310 1.215 6.480 1.375 ;
        RECT  4.840 2.235 6.340 2.395 ;
        RECT  6.150 0.820 6.310 1.375 ;
        RECT  4.465 0.820 6.150 0.980 ;
        RECT  5.570 1.555 5.830 2.050 ;
        RECT  5.420 0.325 5.680 0.595 ;
        RECT  5.220 1.555 5.570 1.715 ;
        RECT  4.555 0.435 5.420 0.595 ;
        RECT  5.060 1.195 5.220 1.715 ;
        RECT  4.960 1.195 5.060 1.355 ;
        RECT  4.580 2.235 4.840 2.560 ;
        RECT  1.665 2.400 4.580 2.560 ;
        RECT  4.395 0.380 4.555 0.595 ;
        RECT  4.305 0.820 4.465 1.950 ;
        RECT  3.870 0.380 4.395 0.540 ;
        RECT  4.210 0.820 4.305 0.980 ;
        RECT  4.050 0.720 4.210 0.980 ;
        RECT  3.815 0.380 3.870 0.910 ;
        RECT  3.710 0.380 3.815 2.100 ;
        RECT  3.655 0.750 3.710 2.100 ;
        RECT  3.455 0.750 3.655 1.010 ;
        RECT  3.145 1.940 3.655 2.100 ;
        RECT  3.275 0.310 3.530 0.470 ;
        RECT  3.115 0.310 3.275 0.810 ;
        RECT  2.885 1.940 3.145 2.220 ;
        RECT  2.635 0.650 3.115 0.810 ;
        RECT  0.695 0.310 2.935 0.470 ;
        RECT  2.095 2.060 2.885 2.220 ;
        RECT  2.475 0.650 2.635 1.880 ;
        RECT  1.625 0.650 2.475 0.810 ;
        RECT  2.375 1.720 2.475 1.880 ;
        RECT  1.935 1.110 2.095 2.220 ;
        RECT  1.485 1.110 1.935 1.270 ;
        RECT  1.405 2.170 1.665 2.560 ;
        RECT  1.150 2.170 1.405 2.330 ;
        RECT  1.150 0.735 1.305 0.995 ;
        RECT  0.990 0.735 1.150 2.330 ;
        RECT  0.535 0.310 0.695 2.180 ;
        RECT  0.125 0.750 0.535 1.010 ;
        RECT  0.385 2.020 0.535 2.180 ;
        RECT  0.125 2.020 0.385 2.280 ;
    END
END DFFHX8MTH

MACRO DFFNHX1MTH
    CLASS CORE ;
    FOREIGN DFFNHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.760 0.765 10.970 1.980 ;
        RECT  10.685 0.765 10.760 1.025 ;
        RECT  10.685 1.720 10.760 1.980 ;
        END
        AntennaDiffArea 0.226 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.905 1.290 10.150 1.580 ;
        RECT  9.745 0.735 9.905 1.990 ;
        RECT  9.585 0.735 9.745 0.995 ;
        END
        AntennaDiffArea 0.26 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.625 1.330 2.235 1.540 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.210 0.425 1.680 ;
        END
        AntennaGateArea 0.1378 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.355 -0.130 11.070 0.130 ;
        RECT  10.095 -0.130 10.355 0.995 ;
        RECT  8.745 -0.130 10.095 0.130 ;
        RECT  8.485 -0.130 8.745 0.300 ;
        RECT  6.885 -0.130 8.485 0.130 ;
        RECT  6.625 -0.130 6.885 0.300 ;
        RECT  5.625 -0.130 6.625 0.130 ;
        RECT  5.365 -0.130 5.625 0.255 ;
        RECT  1.525 -0.130 5.365 0.130 ;
        RECT  0.925 -0.130 1.525 0.415 ;
        RECT  0.000 -0.130 0.925 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.500 2.740 11.070 3.000 ;
        RECT  10.240 2.540 10.500 3.000 ;
        RECT  9.225 2.740 10.240 3.000 ;
        RECT  9.065 1.795 9.225 3.000 ;
        RECT  6.600 2.740 9.065 3.000 ;
        RECT  6.340 2.620 6.600 3.000 ;
        RECT  4.435 2.740 6.340 3.000 ;
        RECT  4.175 2.215 4.435 3.000 ;
        RECT  1.895 2.740 4.175 3.000 ;
        RECT  1.735 2.520 1.895 3.000 ;
        RECT  0.815 2.740 1.735 3.000 ;
        RECT  0.555 2.380 0.815 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.490 1.245 10.580 1.505 ;
        RECT  10.330 1.245 10.490 2.360 ;
        RECT  9.930 2.200 10.330 2.360 ;
        RECT  9.670 2.200 9.930 2.455 ;
        RECT  9.565 2.200 9.670 2.360 ;
        RECT  9.405 1.365 9.565 2.360 ;
        RECT  9.335 1.365 9.405 1.525 ;
        RECT  9.175 0.480 9.335 1.525 ;
        RECT  9.075 0.480 9.175 0.740 ;
        RECT  8.795 1.265 9.175 1.525 ;
        RECT  8.365 0.480 8.525 1.740 ;
        RECT  7.725 0.480 8.365 0.640 ;
        RECT  7.805 0.820 7.965 2.560 ;
        RECT  7.635 0.820 7.805 0.980 ;
        RECT  7.465 0.320 7.725 0.640 ;
        RECT  7.465 1.460 7.625 2.480 ;
        RECT  6.195 0.480 7.465 0.640 ;
        RECT  6.940 2.320 7.465 2.480 ;
        RECT  7.285 0.820 7.385 0.980 ;
        RECT  7.125 0.820 7.285 2.100 ;
        RECT  6.390 1.940 7.125 2.100 ;
        RECT  6.785 0.850 6.945 1.560 ;
        RECT  6.780 2.280 6.940 2.480 ;
        RECT  5.320 0.850 6.785 1.010 ;
        RECT  6.105 2.280 6.780 2.440 ;
        RECT  6.130 1.460 6.390 2.100 ;
        RECT  5.935 0.435 6.195 0.640 ;
        RECT  5.945 2.280 6.105 2.560 ;
        RECT  4.980 2.400 5.945 2.560 ;
        RECT  4.335 0.435 5.935 0.595 ;
        RECT  5.320 1.875 5.660 2.135 ;
        RECT  5.160 0.775 5.320 2.135 ;
        RECT  4.515 0.775 5.160 0.935 ;
        RECT  4.820 1.115 4.980 2.560 ;
        RECT  4.235 1.115 4.820 1.275 ;
        RECT  3.875 1.875 4.820 2.035 ;
        RECT  3.795 1.535 4.635 1.695 ;
        RECT  4.175 0.435 4.335 0.810 ;
        RECT  3.975 0.990 4.235 1.275 ;
        RECT  3.795 0.650 4.175 0.810 ;
        RECT  3.455 0.310 3.995 0.470 ;
        RECT  3.715 1.875 3.875 2.560 ;
        RECT  3.635 0.650 3.795 1.695 ;
        RECT  2.235 2.400 3.715 2.560 ;
        RECT  3.255 1.535 3.635 1.695 ;
        RECT  3.295 0.310 3.455 0.810 ;
        RECT  2.915 0.650 3.295 0.810 ;
        RECT  3.095 1.535 3.255 2.220 ;
        RECT  1.885 0.310 3.115 0.470 ;
        RECT  2.575 2.060 3.095 2.220 ;
        RECT  2.755 0.650 2.915 1.880 ;
        RECT  2.065 0.650 2.755 0.810 ;
        RECT  2.415 0.990 2.575 2.220 ;
        RECT  1.385 0.990 2.415 1.150 ;
        RECT  2.075 1.720 2.235 2.560 ;
        RECT  1.445 1.720 2.075 1.880 ;
        RECT  1.725 0.310 1.885 0.755 ;
        RECT  0.765 0.595 1.725 0.755 ;
        RECT  1.105 2.060 1.665 2.220 ;
        RECT  1.285 1.490 1.445 1.880 ;
        RECT  1.105 0.935 1.385 1.150 ;
        RECT  0.945 0.935 1.105 2.220 ;
        RECT  0.605 0.595 0.765 2.050 ;
        RECT  0.125 0.765 0.605 1.025 ;
        RECT  0.385 1.890 0.605 2.050 ;
        RECT  0.125 1.890 0.385 2.150 ;
    END
END DFFNHX1MTH

MACRO DFFNHX2MTH
    CLASS CORE ;
    FOREIGN DFFNHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.220 0.765 11.380 1.990 ;
        RECT  11.095 0.765 11.220 1.025 ;
        RECT  11.095 1.700 11.220 1.990 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.365 1.290 10.560 1.580 ;
        RECT  10.205 0.380 10.365 1.985 ;
        RECT  10.075 0.380 10.205 0.980 ;
        END
        AntennaDiffArea 0.437 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.330 2.250 1.590 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.475 1.675 ;
        END
        AntennaGateArea 0.1378 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.215 -0.130 11.480 0.130 ;
        RECT  10.615 -0.130 11.215 0.300 ;
        RECT  9.250 -0.130 10.615 0.130 ;
        RECT  8.680 -0.130 9.250 0.300 ;
        RECT  7.190 -0.130 8.680 0.130 ;
        RECT  6.930 -0.130 7.190 0.300 ;
        RECT  6.020 -0.130 6.930 0.130 ;
        RECT  5.760 -0.130 6.020 0.250 ;
        RECT  1.735 -0.130 5.760 0.130 ;
        RECT  0.795 -0.130 1.735 0.275 ;
        RECT  0.000 -0.130 0.795 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.955 2.740 11.480 3.000 ;
        RECT  10.695 2.505 10.955 3.000 ;
        RECT  9.685 2.740 10.695 3.000 ;
        RECT  9.525 1.795 9.685 3.000 ;
        RECT  7.425 2.740 9.525 3.000 ;
        RECT  6.825 2.595 7.425 3.000 ;
        RECT  4.705 2.740 6.825 3.000 ;
        RECT  4.445 2.280 4.705 3.000 ;
        RECT  0.845 2.740 4.445 3.000 ;
        RECT  0.585 2.490 0.845 3.000 ;
        RECT  0.000 2.740 0.585 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.905 1.250 11.030 1.510 ;
        RECT  10.745 1.250 10.905 2.325 ;
        RECT  10.335 2.165 10.745 2.325 ;
        RECT  10.075 2.165 10.335 2.525 ;
        RECT  10.025 2.165 10.075 2.325 ;
        RECT  9.865 1.415 10.025 2.325 ;
        RECT  9.725 1.415 9.865 1.580 ;
        RECT  9.725 0.530 9.825 0.690 ;
        RECT  9.565 0.530 9.725 1.580 ;
        RECT  9.265 1.320 9.565 1.580 ;
        RECT  8.835 0.480 8.995 1.740 ;
        RECT  8.500 0.480 8.835 0.640 ;
        RECT  8.650 2.400 8.750 2.560 ;
        RECT  8.490 0.820 8.650 2.560 ;
        RECT  8.240 0.310 8.500 0.640 ;
        RECT  7.980 0.820 8.490 0.980 ;
        RECT  8.145 1.415 8.305 2.410 ;
        RECT  6.590 0.480 8.240 0.640 ;
        RECT  8.080 1.415 8.145 1.675 ;
        RECT  6.490 2.250 8.145 2.410 ;
        RECT  7.730 1.910 7.965 2.070 ;
        RECT  7.570 0.820 7.730 2.070 ;
        RECT  7.470 0.820 7.570 0.980 ;
        RECT  6.830 1.910 7.570 2.070 ;
        RECT  7.220 1.360 7.390 1.620 ;
        RECT  7.060 0.850 7.220 1.620 ;
        RECT  6.150 0.850 7.060 1.010 ;
        RECT  6.570 1.465 6.830 2.070 ;
        RECT  6.330 0.435 6.590 0.640 ;
        RECT  6.330 2.250 6.490 2.455 ;
        RECT  4.780 0.435 6.330 0.595 ;
        RECT  5.370 2.295 6.330 2.455 ;
        RECT  5.990 0.775 6.150 2.110 ;
        RECT  5.120 0.775 5.990 0.935 ;
        RECT  5.550 1.850 5.990 2.110 ;
        RECT  5.210 1.215 5.370 2.455 ;
        RECT  4.600 1.215 5.210 1.375 ;
        RECT  3.990 1.940 5.210 2.100 ;
        RECT  4.960 0.775 5.120 1.035 ;
        RECT  4.090 1.555 5.030 1.715 ;
        RECT  4.620 0.435 4.780 0.810 ;
        RECT  4.090 0.650 4.620 0.810 ;
        RECT  4.340 0.990 4.600 1.375 ;
        RECT  3.750 0.310 4.440 0.470 ;
        RECT  3.930 0.650 4.090 1.715 ;
        RECT  3.830 1.940 3.990 2.560 ;
        RECT  3.490 1.555 3.930 1.715 ;
        RECT  2.250 2.400 3.830 2.560 ;
        RECT  3.590 0.310 3.750 0.810 ;
        RECT  2.930 0.650 3.590 0.810 ;
        RECT  3.330 1.555 3.490 2.220 ;
        RECT  2.080 0.310 3.410 0.470 ;
        RECT  2.590 2.060 3.330 2.220 ;
        RECT  2.930 1.720 3.030 1.880 ;
        RECT  2.770 0.650 2.930 1.880 ;
        RECT  2.260 0.650 2.770 0.810 ;
        RECT  2.430 0.990 2.590 2.220 ;
        RECT  1.490 0.990 2.430 1.150 ;
        RECT  2.090 1.770 2.250 2.560 ;
        RECT  1.495 1.770 2.090 1.930 ;
        RECT  1.920 0.310 2.080 0.615 ;
        RECT  0.815 0.455 1.920 0.615 ;
        RECT  1.155 2.110 1.695 2.370 ;
        RECT  1.335 1.620 1.495 1.930 ;
        RECT  1.230 0.800 1.490 1.150 ;
        RECT  1.155 0.990 1.230 1.150 ;
        RECT  0.995 0.990 1.155 2.370 ;
        RECT  0.655 0.455 0.815 2.170 ;
        RECT  0.125 0.750 0.655 1.010 ;
        RECT  0.385 2.010 0.655 2.170 ;
        RECT  0.125 2.010 0.385 2.270 ;
    END
END DFFNHX2MTH

MACRO DFFNHX4MTH
    CLASS CORE ;
    FOREIGN DFFNHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.040 0.765 14.250 1.980 ;
        RECT  13.965 0.765 14.040 1.025 ;
        RECT  14.015 1.720 14.040 1.980 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.135 1.685 13.205 1.945 ;
        RECT  12.875 0.385 13.135 1.945 ;
        RECT  12.360 1.290 12.875 1.580 ;
        RECT  12.070 1.290 12.360 1.945 ;
        END
        AntennaDiffArea 0.762 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.450 1.160 2.810 1.540 ;
        END
        AntennaGateArea 0.156 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 1.240 0.720 1.710 ;
        END
        AntennaGateArea 0.1703 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.645 -0.130 14.350 0.130 ;
        RECT  13.385 -0.130 13.645 0.990 ;
        RECT  12.595 -0.130 13.385 0.130 ;
        RECT  12.335 -0.130 12.595 0.525 ;
        RECT  11.640 -0.130 12.335 0.130 ;
        RECT  11.380 -0.130 11.640 0.595 ;
        RECT  7.870 -0.130 11.380 0.130 ;
        RECT  7.610 -0.130 7.870 0.300 ;
        RECT  6.030 -0.130 7.610 0.130 ;
        RECT  5.770 -0.130 6.030 0.975 ;
        RECT  1.785 -0.130 5.770 0.130 ;
        RECT  0.845 -0.130 1.785 0.330 ;
        RECT  0.000 -0.130 0.845 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.745 2.740 14.350 3.000 ;
        RECT  13.485 2.465 13.745 3.000 ;
        RECT  11.550 2.740 13.485 3.000 ;
        RECT  11.390 1.865 11.550 3.000 ;
        RECT  6.720 2.740 11.390 3.000 ;
        RECT  6.460 2.585 6.720 3.000 ;
        RECT  4.610 2.740 6.460 3.000 ;
        RECT  4.350 2.220 4.610 3.000 ;
        RECT  0.740 2.740 4.350 3.000 ;
        RECT  0.570 2.460 0.740 3.000 ;
        RECT  0.000 2.740 0.570 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.675 1.265 13.835 2.285 ;
        RECT  12.210 2.125 13.675 2.285 ;
        RECT  11.890 0.815 12.210 0.975 ;
        RECT  11.950 2.125 12.210 2.540 ;
        RECT  11.890 2.125 11.950 2.285 ;
        RECT  11.730 0.815 11.890 2.285 ;
        RECT  11.320 1.220 11.730 1.480 ;
        RECT  10.980 0.310 11.140 1.735 ;
        RECT  8.930 0.310 10.980 0.470 ;
        RECT  10.700 1.475 10.980 1.735 ;
        RECT  10.640 0.765 10.800 1.280 ;
        RECT  10.220 1.915 10.710 2.075 ;
        RECT  10.220 1.120 10.640 1.280 ;
        RECT  10.080 0.650 10.340 0.940 ;
        RECT  10.060 1.120 10.220 2.480 ;
        RECT  9.275 0.650 10.080 0.810 ;
        RECT  9.830 1.120 10.060 1.280 ;
        RECT  8.950 2.320 10.060 2.480 ;
        RECT  9.570 0.990 9.830 1.280 ;
        RECT  9.275 1.980 9.510 2.140 ;
        RECT  9.115 0.650 9.275 2.140 ;
        RECT  9.110 0.650 9.115 1.275 ;
        RECT  8.410 1.115 9.110 1.275 ;
        RECT  8.790 2.220 8.950 2.480 ;
        RECT  8.770 0.310 8.930 0.640 ;
        RECT  7.180 0.480 8.770 0.640 ;
        RECT  8.450 1.455 8.610 2.475 ;
        RECT  7.790 2.315 8.450 2.475 ;
        RECT  8.270 0.820 8.410 1.275 ;
        RECT  8.110 0.820 8.270 2.135 ;
        RECT  7.970 1.905 8.110 2.135 ;
        RECT  7.070 1.905 7.970 2.065 ;
        RECT  7.770 0.865 7.930 1.525 ;
        RECT  7.630 2.245 7.790 2.475 ;
        RECT  6.710 0.865 7.770 1.025 ;
        RECT  6.175 2.245 7.630 2.405 ;
        RECT  6.920 0.345 7.180 0.640 ;
        RECT  6.910 1.340 7.070 2.065 ;
        RECT  6.370 0.480 6.920 0.640 ;
        RECT  6.550 0.865 6.710 1.655 ;
        RECT  5.930 1.495 6.550 1.655 ;
        RECT  6.210 0.480 6.370 1.315 ;
        RECT  5.550 1.155 6.210 1.315 ;
        RECT  6.015 2.245 6.175 2.445 ;
        RECT  4.975 2.285 6.015 2.445 ;
        RECT  5.330 1.495 5.930 2.085 ;
        RECT  5.390 0.465 5.550 1.315 ;
        RECT  4.640 0.465 5.390 0.625 ;
        RECT  5.210 1.495 5.330 1.655 ;
        RECT  5.050 0.805 5.210 1.655 ;
        RECT  4.820 0.805 5.050 0.965 ;
        RECT  4.870 1.880 4.975 2.445 ;
        RECT  4.815 1.145 4.870 2.445 ;
        RECT  4.710 1.145 4.815 2.040 ;
        RECT  4.465 1.145 4.710 1.305 ;
        RECT  3.830 1.880 4.710 2.040 ;
        RECT  4.480 0.465 4.640 0.810 ;
        RECT  4.025 1.540 4.530 1.700 ;
        RECT  4.025 0.650 4.480 0.810 ;
        RECT  4.205 0.990 4.465 1.305 ;
        RECT  3.685 0.310 4.300 0.470 ;
        RECT  3.865 0.650 4.025 1.700 ;
        RECT  3.490 1.540 3.865 1.700 ;
        RECT  3.670 1.880 3.830 2.560 ;
        RECT  3.525 0.310 3.685 0.810 ;
        RECT  1.930 2.400 3.670 2.560 ;
        RECT  3.150 0.650 3.525 0.810 ;
        RECT  3.330 1.540 3.490 2.220 ;
        RECT  2.125 0.310 3.345 0.470 ;
        RECT  2.270 2.060 3.330 2.220 ;
        RECT  2.990 0.650 3.150 1.880 ;
        RECT  2.305 0.650 2.990 0.810 ;
        RECT  2.565 1.720 2.990 1.880 ;
        RECT  2.110 0.990 2.270 2.220 ;
        RECT  1.965 0.310 2.125 0.810 ;
        RECT  1.585 0.990 2.110 1.150 ;
        RECT  1.120 0.650 1.965 0.810 ;
        RECT  1.770 1.540 1.930 2.560 ;
        RECT  1.425 0.990 1.585 2.265 ;
        RECT  1.300 0.990 1.425 1.250 ;
        RECT  0.960 0.650 1.120 2.070 ;
        RECT  0.165 0.765 0.960 1.025 ;
        RECT  0.385 1.910 0.960 2.070 ;
        RECT  0.125 1.910 0.385 2.170 ;
    END
END DFFNHX4MTH

MACRO DFFNHX8MTH
    CLASS CORE ;
    FOREIGN DFFNHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.270 0.765 15.480 1.980 ;
        RECT  15.185 0.765 15.270 1.025 ;
        RECT  15.195 1.720 15.270 1.980 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.105 0.385 14.365 1.945 ;
        RECT  13.345 1.290 14.105 1.580 ;
        RECT  13.285 0.385 13.345 1.580 ;
        RECT  13.085 0.385 13.285 1.945 ;
        RECT  13.025 1.290 13.085 1.945 ;
        RECT  12.360 1.290 13.025 1.580 ;
        RECT  12.070 1.290 12.360 1.945 ;
        END
        AntennaDiffArea 1.362 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.450 1.160 2.810 1.540 ;
        END
        AntennaGateArea 0.2912 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 1.240 0.720 1.710 ;
        END
        AntennaGateArea 0.273 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.875 -0.130 15.580 0.130 ;
        RECT  14.615 -0.130 14.875 0.985 ;
        RECT  13.855 -0.130 14.615 0.130 ;
        RECT  13.595 -0.130 13.855 0.985 ;
        RECT  12.835 -0.130 13.595 0.130 ;
        RECT  12.575 -0.130 12.835 0.985 ;
        RECT  11.740 -0.130 12.575 0.130 ;
        RECT  11.480 -0.130 11.740 0.635 ;
        RECT  7.870 -0.130 11.480 0.130 ;
        RECT  7.610 -0.130 7.870 0.300 ;
        RECT  6.030 -0.130 7.610 0.130 ;
        RECT  5.770 -0.130 6.030 0.975 ;
        RECT  1.720 -0.130 5.770 0.130 ;
        RECT  0.780 -0.130 1.720 0.330 ;
        RECT  0.000 -0.130 0.780 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.915 2.740 15.580 3.000 ;
        RECT  14.655 2.465 14.915 3.000 ;
        RECT  13.825 2.740 14.655 3.000 ;
        RECT  13.565 2.465 13.825 3.000 ;
        RECT  12.775 2.740 13.565 3.000 ;
        RECT  12.515 2.465 12.775 3.000 ;
        RECT  11.550 2.740 12.515 3.000 ;
        RECT  11.390 1.895 11.550 3.000 ;
        RECT  6.720 2.740 11.390 3.000 ;
        RECT  6.460 2.585 6.720 3.000 ;
        RECT  4.610 2.740 6.460 3.000 ;
        RECT  4.350 2.220 4.610 3.000 ;
        RECT  0.000 2.740 4.350 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.920 1.225 15.090 1.485 ;
        RECT  14.760 1.225 14.920 2.285 ;
        RECT  12.210 2.125 14.760 2.285 ;
        RECT  11.890 0.815 12.315 0.975 ;
        RECT  11.950 2.125 12.210 2.540 ;
        RECT  11.890 2.125 11.950 2.285 ;
        RECT  11.730 0.815 11.890 2.285 ;
        RECT  11.320 1.220 11.730 1.480 ;
        RECT  10.980 0.310 11.140 1.735 ;
        RECT  8.930 0.310 10.980 0.470 ;
        RECT  10.700 1.475 10.980 1.735 ;
        RECT  10.640 0.765 10.800 1.280 ;
        RECT  10.220 1.945 10.710 2.105 ;
        RECT  10.220 1.120 10.640 1.280 ;
        RECT  10.220 2.400 10.600 2.560 ;
        RECT  10.080 0.650 10.340 0.940 ;
        RECT  10.060 1.120 10.220 2.560 ;
        RECT  9.290 0.650 10.080 0.810 ;
        RECT  9.830 1.120 10.060 1.280 ;
        RECT  8.950 2.400 10.060 2.560 ;
        RECT  9.570 0.990 9.830 1.280 ;
        RECT  9.290 1.980 9.510 2.140 ;
        RECT  9.130 0.650 9.290 2.140 ;
        RECT  9.110 0.650 9.130 1.275 ;
        RECT  8.410 1.115 9.110 1.275 ;
        RECT  8.790 1.880 8.950 2.560 ;
        RECT  8.770 0.310 8.930 0.640 ;
        RECT  7.180 0.480 8.770 0.640 ;
        RECT  8.450 1.480 8.610 2.475 ;
        RECT  7.790 2.315 8.450 2.475 ;
        RECT  8.270 0.820 8.410 1.275 ;
        RECT  8.110 0.820 8.270 2.135 ;
        RECT  7.970 1.905 8.110 2.135 ;
        RECT  7.070 1.905 7.970 2.065 ;
        RECT  7.770 0.865 7.930 1.525 ;
        RECT  7.630 2.245 7.790 2.475 ;
        RECT  6.710 0.865 7.770 1.025 ;
        RECT  6.175 2.245 7.630 2.405 ;
        RECT  6.920 0.310 7.180 0.640 ;
        RECT  6.910 1.340 7.070 2.065 ;
        RECT  6.370 0.480 6.920 0.640 ;
        RECT  6.550 0.865 6.710 1.655 ;
        RECT  5.930 1.495 6.550 1.655 ;
        RECT  6.210 0.480 6.370 1.315 ;
        RECT  5.550 1.155 6.210 1.315 ;
        RECT  6.015 2.245 6.175 2.455 ;
        RECT  4.975 2.295 6.015 2.455 ;
        RECT  5.330 1.495 5.930 2.085 ;
        RECT  5.390 0.465 5.550 1.315 ;
        RECT  4.640 0.465 5.390 0.625 ;
        RECT  5.210 1.495 5.330 1.655 ;
        RECT  5.050 0.805 5.210 1.655 ;
        RECT  4.820 0.805 5.050 0.965 ;
        RECT  4.870 1.880 4.975 2.455 ;
        RECT  4.815 1.145 4.870 2.455 ;
        RECT  4.710 1.145 4.815 2.040 ;
        RECT  4.465 1.145 4.710 1.305 ;
        RECT  3.830 1.880 4.710 2.040 ;
        RECT  4.480 0.465 4.640 0.810 ;
        RECT  4.025 1.540 4.530 1.700 ;
        RECT  4.025 0.650 4.480 0.810 ;
        RECT  4.205 0.990 4.465 1.305 ;
        RECT  3.685 0.310 4.300 0.470 ;
        RECT  3.865 0.650 4.025 1.700 ;
        RECT  3.490 1.540 3.865 1.700 ;
        RECT  3.670 1.880 3.830 2.560 ;
        RECT  3.525 0.310 3.685 0.810 ;
        RECT  1.930 2.400 3.670 2.560 ;
        RECT  3.150 0.650 3.525 0.810 ;
        RECT  3.330 1.540 3.490 2.220 ;
        RECT  2.060 0.310 3.345 0.470 ;
        RECT  2.270 2.060 3.330 2.220 ;
        RECT  2.990 0.650 3.150 1.880 ;
        RECT  2.240 0.650 2.990 0.810 ;
        RECT  2.565 1.720 2.990 1.880 ;
        RECT  2.110 0.990 2.270 2.220 ;
        RECT  1.585 0.990 2.110 1.150 ;
        RECT  1.900 0.310 2.060 0.810 ;
        RECT  1.770 1.540 1.930 2.560 ;
        RECT  1.120 0.650 1.900 0.810 ;
        RECT  1.425 0.990 1.585 2.515 ;
        RECT  1.300 0.990 1.425 1.250 ;
        RECT  0.960 0.650 1.120 2.180 ;
        RECT  0.425 0.650 0.960 0.810 ;
        RECT  0.385 2.020 0.960 2.180 ;
        RECT  0.165 0.650 0.425 0.910 ;
        RECT  0.125 2.020 0.385 2.280 ;
    END
END DFFNHX8MTH

MACRO DFFNSRHX1MTH
    CLASS CORE ;
    FOREIGN DFFNSRHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.145 4.065 1.660 ;
        END
        AntennaGateArea 0.1391 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 1.385 10.445 1.545 ;
        RECT  8.880 1.385 9.040 1.635 ;
        RECT  8.140 1.475 8.880 1.635 ;
        RECT  7.440 1.330 8.140 1.635 ;
        END
        AntennaGateArea 0.1417 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.365 2.255 13.095 2.415 ;
        RECT  12.365 0.815 12.650 1.130 ;
        RECT  12.205 0.815 12.365 2.415 ;
        END
        AntennaDiffArea 0.348 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.015 0.740 14.250 2.285 ;
        END
        AntennaDiffArea 0.34 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.385 1.255 2.675 1.520 ;
        RECT  2.145 1.255 2.385 1.990 ;
        END
        AntennaGateArea 0.0676 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.240 1.015 1.580 ;
        END
        AntennaGateArea 0.1469 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.525 -0.130 14.350 0.130 ;
        RECT  12.925 -0.130 13.525 0.260 ;
        RECT  2.360 -0.130 12.925 0.130 ;
        RECT  1.760 -0.130 2.360 0.250 ;
        RECT  0.810 -0.130 1.760 0.130 ;
        RECT  0.210 -0.130 0.810 0.250 ;
        RECT  0.000 -0.130 0.210 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.715 2.740 14.350 3.000 ;
        RECT  13.455 1.685 13.715 3.000 ;
        RECT  8.230 2.740 13.455 3.000 ;
        RECT  7.970 2.620 8.230 3.000 ;
        RECT  7.290 2.740 7.970 3.000 ;
        RECT  7.030 2.620 7.290 3.000 ;
        RECT  6.140 2.740 7.030 3.000 ;
        RECT  5.880 2.620 6.140 3.000 ;
        RECT  5.285 2.740 5.880 3.000 ;
        RECT  5.025 2.620 5.285 3.000 ;
        RECT  2.565 2.740 5.025 3.000 ;
        RECT  2.405 2.530 2.565 3.000 ;
        RECT  0.755 2.740 2.405 3.000 ;
        RECT  0.255 2.365 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.665 1.185 13.825 1.445 ;
        RECT  13.505 0.475 13.665 1.445 ;
        RECT  12.000 0.475 13.505 0.635 ;
        RECT  13.325 1.185 13.505 1.445 ;
        RECT  13.095 0.815 13.185 0.975 ;
        RECT  12.925 0.815 13.095 1.945 ;
        RECT  12.545 1.310 12.925 1.945 ;
        RECT  11.840 0.355 12.000 2.505 ;
        RECT  11.435 0.355 11.840 0.550 ;
        RECT  11.240 2.295 11.840 2.505 ;
        RECT  11.500 0.760 11.660 2.115 ;
        RECT  11.360 0.760 11.500 0.920 ;
        RECT  10.785 1.955 11.500 2.115 ;
        RECT  9.560 0.355 11.435 0.515 ;
        RECT  9.950 2.295 11.240 2.455 ;
        RECT  11.020 0.695 11.180 1.775 ;
        RECT  9.380 0.695 11.020 0.855 ;
        RECT  10.625 1.035 10.785 2.115 ;
        RECT  9.040 1.035 10.625 1.195 ;
        RECT  10.180 1.865 10.625 2.115 ;
        RECT  8.910 1.815 9.670 1.975 ;
        RECT  9.125 2.185 9.385 2.440 ;
        RECT  9.220 0.310 9.380 0.855 ;
        RECT  2.710 0.310 9.220 0.470 ;
        RECT  6.700 2.280 9.125 2.440 ;
        RECT  8.880 0.650 9.040 1.195 ;
        RECT  8.750 1.815 8.910 2.100 ;
        RECT  3.610 0.650 8.880 0.810 ;
        RECT  7.130 1.940 8.750 2.100 ;
        RECT  8.540 0.990 8.700 1.250 ;
        RECT  7.130 0.990 8.540 1.150 ;
        RECT  6.970 0.990 7.130 2.100 ;
        RECT  6.440 2.280 6.700 2.560 ;
        RECT  6.530 1.075 6.690 2.100 ;
        RECT  5.740 1.940 6.530 2.100 ;
        RECT  4.845 2.280 6.440 2.440 ;
        RECT  5.580 0.990 5.740 2.100 ;
        RECT  5.390 0.990 5.580 1.150 ;
        RECT  5.280 1.940 5.580 2.100 ;
        RECT  5.210 1.335 5.400 1.595 ;
        RECT  5.020 1.910 5.280 2.100 ;
        RECT  5.050 1.130 5.210 1.595 ;
        RECT  4.500 1.130 5.050 1.290 ;
        RECT  4.840 1.470 4.870 1.730 ;
        RECT  4.840 2.280 4.845 2.555 ;
        RECT  4.680 1.470 4.840 2.555 ;
        RECT  2.905 2.395 4.680 2.555 ;
        RECT  4.340 1.130 4.500 2.215 ;
        RECT  3.270 2.055 4.340 2.215 ;
        RECT  3.450 0.650 3.610 1.875 ;
        RECT  3.400 0.650 3.450 0.810 ;
        RECT  3.150 1.665 3.270 2.215 ;
        RECT  3.110 0.650 3.150 2.215 ;
        RECT  2.990 0.650 3.110 1.895 ;
        RECT  2.890 0.650 2.990 0.810 ;
        RECT  2.890 1.735 2.990 1.895 ;
        RECT  2.745 2.180 2.905 2.555 ;
        RECT  2.110 2.180 2.745 2.345 ;
        RECT  2.550 0.310 2.710 0.590 ;
        RECT  1.605 0.430 2.550 0.590 ;
        RECT  1.965 2.180 2.110 2.485 ;
        RECT  1.965 0.815 2.075 0.975 ;
        RECT  1.785 0.815 1.965 2.485 ;
        RECT  1.625 1.285 1.785 1.545 ;
        RECT  1.445 0.430 1.605 1.010 ;
        RECT  1.415 1.740 1.605 2.000 ;
        RECT  1.415 0.850 1.445 1.010 ;
        RECT  1.195 0.850 1.415 2.000 ;
        RECT  1.005 0.310 1.265 0.670 ;
        RECT  0.385 0.490 1.005 0.670 ;
        RECT  0.330 0.490 0.385 1.025 ;
        RECT  0.330 1.740 0.365 2.000 ;
        RECT  0.125 0.490 0.330 2.000 ;
    END
END DFFNSRHX1MTH

MACRO DFFNSRHX2MTH
    CLASS CORE ;
    FOREIGN DFFNSRHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.145 4.065 1.660 ;
        END
        AntennaGateArea 0.1612 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 1.385 10.445 1.545 ;
        RECT  8.880 1.385 9.040 1.635 ;
        RECT  8.140 1.475 8.880 1.635 ;
        RECT  7.710 1.330 8.140 1.635 ;
        END
        AntennaGateArea 0.1716 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.610 2.255 13.095 2.415 ;
        RECT  12.365 2.065 12.610 2.415 ;
        RECT  12.365 0.815 12.465 0.975 ;
        RECT  12.205 0.815 12.365 2.415 ;
        END
        AntennaDiffArea 0.348 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.015 0.400 14.250 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.255 2.675 1.580 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.225 0.895 1.580 ;
        END
        AntennaGateArea 0.1469 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.520 -0.130 14.350 0.130 ;
        RECT  12.920 -0.130 13.520 0.260 ;
        RECT  2.370 -0.130 12.920 0.130 ;
        RECT  1.770 -0.130 2.370 0.250 ;
        RECT  0.810 -0.130 1.770 0.130 ;
        RECT  0.210 -0.130 0.810 0.250 ;
        RECT  0.000 -0.130 0.210 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.715 2.740 14.350 3.000 ;
        RECT  13.455 1.830 13.715 3.000 ;
        RECT  8.230 2.740 13.455 3.000 ;
        RECT  7.970 2.620 8.230 3.000 ;
        RECT  7.290 2.740 7.970 3.000 ;
        RECT  7.030 2.620 7.290 3.000 ;
        RECT  6.140 2.740 7.030 3.000 ;
        RECT  5.880 2.620 6.140 3.000 ;
        RECT  5.285 2.740 5.880 3.000 ;
        RECT  5.025 2.620 5.285 3.000 ;
        RECT  2.565 2.740 5.025 3.000 ;
        RECT  2.405 2.530 2.565 3.000 ;
        RECT  0.755 2.740 2.405 3.000 ;
        RECT  0.255 2.365 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.665 1.185 13.825 1.445 ;
        RECT  13.505 0.475 13.665 1.445 ;
        RECT  12.000 0.475 13.505 0.635 ;
        RECT  13.325 1.185 13.505 1.445 ;
        RECT  13.095 0.815 13.195 0.975 ;
        RECT  12.935 0.815 13.095 1.945 ;
        RECT  12.545 1.240 12.935 1.840 ;
        RECT  11.840 0.355 12.000 2.505 ;
        RECT  11.435 0.355 11.840 0.550 ;
        RECT  11.240 2.295 11.840 2.505 ;
        RECT  11.500 0.760 11.660 2.115 ;
        RECT  11.360 0.760 11.500 0.920 ;
        RECT  10.785 1.955 11.500 2.115 ;
        RECT  9.560 0.355 11.435 0.515 ;
        RECT  9.950 2.295 11.240 2.455 ;
        RECT  11.020 0.695 11.180 1.775 ;
        RECT  9.380 0.695 11.020 0.855 ;
        RECT  10.625 1.035 10.785 2.115 ;
        RECT  9.040 1.035 10.625 1.195 ;
        RECT  10.180 1.865 10.625 2.115 ;
        RECT  8.910 1.815 9.670 1.975 ;
        RECT  9.125 2.185 9.385 2.440 ;
        RECT  9.220 0.310 9.380 0.855 ;
        RECT  2.710 0.310 9.220 0.470 ;
        RECT  6.700 2.280 9.125 2.440 ;
        RECT  8.880 0.650 9.040 1.195 ;
        RECT  8.750 1.815 8.910 2.100 ;
        RECT  3.610 0.650 8.880 0.810 ;
        RECT  7.130 1.940 8.750 2.100 ;
        RECT  8.540 0.990 8.700 1.250 ;
        RECT  7.130 0.990 8.540 1.150 ;
        RECT  6.970 0.990 7.130 2.100 ;
        RECT  6.440 2.280 6.700 2.560 ;
        RECT  6.530 1.075 6.690 2.100 ;
        RECT  6.240 1.840 6.530 2.100 ;
        RECT  4.845 2.280 6.440 2.440 ;
        RECT  5.740 1.840 6.240 2.000 ;
        RECT  5.580 0.990 5.740 2.000 ;
        RECT  5.390 0.990 5.580 1.150 ;
        RECT  5.280 1.840 5.580 2.000 ;
        RECT  5.210 1.335 5.400 1.595 ;
        RECT  5.020 1.840 5.280 2.070 ;
        RECT  5.050 1.130 5.210 1.595 ;
        RECT  4.500 1.130 5.050 1.290 ;
        RECT  4.840 1.470 4.870 1.730 ;
        RECT  4.840 2.280 4.845 2.555 ;
        RECT  4.710 1.470 4.840 2.555 ;
        RECT  4.680 1.540 4.710 2.555 ;
        RECT  2.905 2.395 4.680 2.555 ;
        RECT  4.340 1.130 4.500 2.215 ;
        RECT  3.270 2.055 4.340 2.215 ;
        RECT  3.450 0.650 3.610 1.875 ;
        RECT  3.400 0.650 3.450 0.810 ;
        RECT  3.155 1.665 3.270 2.215 ;
        RECT  3.110 0.740 3.155 2.215 ;
        RECT  2.995 0.740 3.110 1.895 ;
        RECT  2.890 0.740 2.995 0.900 ;
        RECT  2.890 1.735 2.995 1.895 ;
        RECT  2.745 2.085 2.905 2.555 ;
        RECT  2.110 2.085 2.745 2.250 ;
        RECT  2.550 0.310 2.710 0.635 ;
        RECT  1.605 0.475 2.550 0.635 ;
        RECT  1.965 2.085 2.110 2.485 ;
        RECT  1.965 0.815 2.075 0.975 ;
        RECT  1.785 0.815 1.965 2.485 ;
        RECT  1.625 1.285 1.785 1.545 ;
        RECT  1.445 0.475 1.605 1.010 ;
        RECT  1.415 1.740 1.605 2.000 ;
        RECT  1.415 0.850 1.445 1.010 ;
        RECT  1.195 0.850 1.415 2.000 ;
        RECT  1.005 0.310 1.265 0.670 ;
        RECT  0.385 0.490 1.005 0.670 ;
        RECT  0.330 0.490 0.385 1.025 ;
        RECT  0.330 1.740 0.365 2.000 ;
        RECT  0.125 0.490 0.330 2.000 ;
    END
END DFFNSRHX2MTH

MACRO DFFNSRHX4MTH
    CLASS CORE ;
    FOREIGN DFFNSRHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.760 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.230 4.140 1.760 ;
        END
        AntennaGateArea 0.1807 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.040 1.385 10.445 1.545 ;
        RECT  8.880 1.385 9.040 1.635 ;
        RECT  8.140 1.475 8.880 1.635 ;
        RECT  7.645 1.330 8.140 1.635 ;
        END
        AntennaGateArea 0.2093 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.610 2.255 13.075 2.415 ;
        RECT  12.345 2.065 12.610 2.415 ;
        RECT  12.345 0.815 12.465 0.975 ;
        RECT  12.185 0.815 12.345 2.415 ;
        END
        AntennaDiffArea 0.384 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.235 1.290 14.325 1.580 ;
        RECT  14.040 0.400 14.235 2.285 ;
        RECT  13.915 0.400 14.040 1.000 ;
        RECT  13.915 1.685 14.040 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.150 2.675 1.410 ;
        RECT  2.145 1.150 2.360 1.990 ;
        END
        AntennaGateArea 0.156 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.225 0.895 1.580 ;
        END
        AntennaGateArea 0.1664 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.585 -0.130 14.760 0.130 ;
        RECT  14.425 -0.130 14.585 1.000 ;
        RECT  13.520 -0.130 14.425 0.130 ;
        RECT  12.920 -0.130 13.520 0.260 ;
        RECT  4.370 -0.130 12.920 0.130 ;
        RECT  4.110 -0.130 4.370 0.250 ;
        RECT  0.785 -0.130 4.110 0.130 ;
        RECT  0.185 -0.130 0.785 0.250 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.585 2.740 14.760 3.000 ;
        RECT  14.425 1.815 14.585 3.000 ;
        RECT  13.585 2.740 14.425 3.000 ;
        RECT  13.325 2.195 13.585 3.000 ;
        RECT  7.005 2.740 13.325 3.000 ;
        RECT  6.745 2.620 7.005 3.000 ;
        RECT  6.065 2.740 6.745 3.000 ;
        RECT  5.805 2.620 6.065 3.000 ;
        RECT  4.185 2.740 5.805 3.000 ;
        RECT  3.585 2.620 4.185 3.000 ;
        RECT  2.615 2.740 3.585 3.000 ;
        RECT  2.355 2.620 2.615 3.000 ;
        RECT  0.755 2.740 2.355 3.000 ;
        RECT  0.255 2.365 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.665 1.185 13.825 1.445 ;
        RECT  13.505 0.475 13.665 1.445 ;
        RECT  12.000 0.475 13.505 0.635 ;
        RECT  13.325 1.185 13.505 1.445 ;
        RECT  12.845 0.815 13.105 1.945 ;
        RECT  12.525 1.240 12.845 1.840 ;
        RECT  11.840 0.355 12.000 2.505 ;
        RECT  11.435 0.355 11.840 0.550 ;
        RECT  11.220 2.295 11.840 2.505 ;
        RECT  11.500 0.760 11.660 2.115 ;
        RECT  11.360 0.760 11.500 0.920 ;
        RECT  10.785 1.955 11.500 2.115 ;
        RECT  9.550 0.355 11.435 0.515 ;
        RECT  9.940 2.295 11.220 2.455 ;
        RECT  11.020 0.695 11.180 1.775 ;
        RECT  9.370 0.695 11.020 0.855 ;
        RECT  10.625 1.035 10.785 2.115 ;
        RECT  9.030 1.035 10.625 1.195 ;
        RECT  10.170 1.865 10.625 2.115 ;
        RECT  8.910 1.815 9.660 1.975 ;
        RECT  9.140 2.185 9.400 2.560 ;
        RECT  9.210 0.310 9.370 0.855 ;
        RECT  4.825 0.310 9.210 0.470 ;
        RECT  7.345 2.400 9.140 2.560 ;
        RECT  8.870 0.650 9.030 1.195 ;
        RECT  8.750 1.815 8.910 2.195 ;
        RECT  5.165 0.650 8.870 0.810 ;
        RECT  7.795 2.035 8.750 2.195 ;
        RECT  8.530 0.990 8.690 1.250 ;
        RECT  7.065 0.990 8.530 1.150 ;
        RECT  7.535 1.940 7.795 2.195 ;
        RECT  7.065 1.940 7.535 2.100 ;
        RECT  7.185 2.280 7.345 2.560 ;
        RECT  6.535 2.280 7.185 2.440 ;
        RECT  6.905 0.990 7.065 2.100 ;
        RECT  6.565 1.025 6.725 2.100 ;
        RECT  6.175 1.860 6.565 2.100 ;
        RECT  6.270 2.280 6.535 2.560 ;
        RECT  5.570 2.280 6.270 2.440 ;
        RECT  5.650 1.860 6.175 2.020 ;
        RECT  5.490 0.990 5.650 2.020 ;
        RECT  5.410 2.280 5.570 2.480 ;
        RECT  5.345 0.990 5.490 1.150 ;
        RECT  5.230 1.860 5.490 2.020 ;
        RECT  4.825 2.320 5.410 2.480 ;
        RECT  5.165 1.335 5.310 1.595 ;
        RECT  5.005 1.860 5.230 2.120 ;
        RECT  5.005 0.650 5.165 0.950 ;
        RECT  5.005 1.130 5.165 1.595 ;
        RECT  3.610 0.790 5.005 0.950 ;
        RECT  4.485 1.130 5.005 1.290 ;
        RECT  4.665 0.310 4.825 0.610 ;
        RECT  4.665 1.485 4.825 2.480 ;
        RECT  3.940 0.450 4.665 0.610 ;
        RECT  2.075 2.280 4.665 2.440 ;
        RECT  4.325 1.130 4.485 2.100 ;
        RECT  3.155 1.940 4.325 2.100 ;
        RECT  3.780 0.310 3.940 0.610 ;
        RECT  1.605 0.310 3.780 0.470 ;
        RECT  3.350 0.680 3.610 1.760 ;
        RECT  2.995 0.650 3.155 2.100 ;
        RECT  2.840 0.650 2.995 0.810 ;
        RECT  2.890 1.690 2.995 2.100 ;
        RECT  1.965 0.650 2.075 0.810 ;
        RECT  1.965 2.280 2.075 2.525 ;
        RECT  1.785 0.650 1.965 2.525 ;
        RECT  1.575 1.285 1.785 1.545 ;
        RECT  1.445 0.310 1.605 1.010 ;
        RECT  1.305 1.740 1.605 2.000 ;
        RECT  1.305 0.790 1.445 1.010 ;
        RECT  1.095 0.790 1.305 2.000 ;
        RECT  1.005 0.310 1.265 0.610 ;
        RECT  0.385 0.430 1.005 0.610 ;
        RECT  0.310 0.430 0.385 1.025 ;
        RECT  0.310 1.740 0.335 2.000 ;
        RECT  0.125 0.430 0.310 2.000 ;
    END
END DFFNSRHX4MTH

MACRO DFFNSRHX8MTH
    CLASS CORE ;
    FOREIGN DFFNSRHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 1.230 4.475 1.740 ;
        END
        AntennaGateArea 0.2249 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.435 1.395 10.840 1.555 ;
        RECT  9.275 1.395 9.435 1.635 ;
        RECT  8.550 1.475 9.275 1.635 ;
        RECT  8.105 1.330 8.550 1.635 ;
        END
        AntennaGateArea 0.2119 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.760 2.150 13.675 2.415 ;
        RECT  12.760 0.815 12.860 0.975 ;
        RECT  12.600 0.815 12.760 2.415 ;
        END
        AntennaDiffArea 0.398 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.455 0.400 15.725 2.285 ;
        RECT  14.695 0.905 15.455 1.065 ;
        RECT  15.025 1.330 15.455 1.745 ;
        RECT  14.695 1.585 15.025 1.745 ;
        RECT  14.435 0.400 14.695 1.065 ;
        RECT  14.435 1.585 14.695 2.285 ;
        END
        AntennaDiffArea 1.204 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 0.990 3.105 1.315 ;
        RECT  2.560 0.990 2.770 1.655 ;
        END
        AntennaGateArea 0.2041 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.195 0.925 1.580 ;
        END
        AntennaGateArea 0.2951 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.225 -0.130 16.400 0.130 ;
        RECT  15.965 -0.130 16.225 1.000 ;
        RECT  15.205 -0.130 15.965 0.130 ;
        RECT  14.945 -0.130 15.205 0.705 ;
        RECT  13.955 -0.130 14.945 0.130 ;
        RECT  13.355 -0.130 13.955 0.260 ;
        RECT  4.750 -0.130 13.355 0.130 ;
        RECT  4.550 -0.130 4.750 0.300 ;
        RECT  0.925 -0.130 4.550 0.130 ;
        RECT  0.665 -0.130 0.925 0.250 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.225 2.740 16.400 3.000 ;
        RECT  15.965 1.815 16.225 3.000 ;
        RECT  15.205 2.740 15.965 3.000 ;
        RECT  14.945 1.925 15.205 3.000 ;
        RECT  14.155 2.740 14.945 3.000 ;
        RECT  13.895 2.230 14.155 3.000 ;
        RECT  11.515 2.740 13.895 3.000 ;
        RECT  11.255 2.620 11.515 3.000 ;
        RECT  7.685 2.740 11.255 3.000 ;
        RECT  7.425 2.620 7.685 3.000 ;
        RECT  6.535 2.740 7.425 3.000 ;
        RECT  6.275 2.620 6.535 3.000 ;
        RECT  4.570 2.740 6.275 3.000 ;
        RECT  3.970 2.620 4.570 3.000 ;
        RECT  1.985 2.740 3.970 3.000 ;
        RECT  1.785 2.255 1.985 3.000 ;
        RECT  0.735 2.740 1.785 3.000 ;
        RECT  0.235 2.530 0.735 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.145 1.245 14.670 1.405 ;
        RECT  13.985 0.475 14.145 1.405 ;
        RECT  12.395 0.475 13.985 0.635 ;
        RECT  13.730 1.245 13.985 1.405 ;
        RECT  13.490 1.685 13.600 1.945 ;
        RECT  13.490 0.815 13.540 0.975 ;
        RECT  13.280 0.815 13.490 1.945 ;
        RECT  12.940 1.240 13.280 1.945 ;
        RECT  12.235 0.355 12.395 2.505 ;
        RECT  11.830 0.355 12.235 0.565 ;
        RECT  11.765 2.280 12.235 2.505 ;
        RECT  11.895 0.775 12.055 2.100 ;
        RECT  11.755 0.775 11.895 0.935 ;
        RECT  11.180 1.940 11.895 2.100 ;
        RECT  9.955 0.355 11.830 0.515 ;
        RECT  10.345 2.280 11.765 2.440 ;
        RECT  11.525 1.600 11.625 1.760 ;
        RECT  11.365 0.695 11.525 1.760 ;
        RECT  9.775 0.695 11.365 0.855 ;
        RECT  11.020 1.035 11.180 2.100 ;
        RECT  9.435 1.035 11.020 1.195 ;
        RECT  10.575 1.865 11.020 2.100 ;
        RECT  9.305 1.815 10.065 1.975 ;
        RECT  9.545 2.185 9.805 2.440 ;
        RECT  9.615 0.310 9.775 0.855 ;
        RECT  5.150 0.310 9.615 0.470 ;
        RECT  7.095 2.280 9.545 2.440 ;
        RECT  9.275 0.650 9.435 1.195 ;
        RECT  9.145 1.815 9.305 2.100 ;
        RECT  5.565 0.650 9.275 0.810 ;
        RECT  7.525 1.940 9.145 2.100 ;
        RECT  8.935 0.990 9.095 1.250 ;
        RECT  7.525 0.990 8.935 1.150 ;
        RECT  7.365 0.990 7.525 2.100 ;
        RECT  7.025 0.990 7.185 2.100 ;
        RECT  6.835 2.280 7.095 2.560 ;
        RECT  6.635 1.860 7.025 2.100 ;
        RECT  5.965 2.280 6.835 2.440 ;
        RECT  6.135 1.860 6.635 2.020 ;
        RECT  5.975 0.990 6.135 2.020 ;
        RECT  5.785 0.990 5.975 1.150 ;
        RECT  5.625 1.860 5.975 2.020 ;
        RECT  5.805 2.280 5.965 2.480 ;
        RECT  5.265 2.320 5.805 2.480 ;
        RECT  5.605 1.335 5.795 1.595 ;
        RECT  5.465 1.860 5.625 2.120 ;
        RECT  5.445 1.160 5.605 1.595 ;
        RECT  5.405 0.650 5.565 0.980 ;
        RECT  4.825 1.160 5.445 1.320 ;
        RECT  4.015 0.820 5.405 0.980 ;
        RECT  5.105 1.535 5.265 2.480 ;
        RECT  4.990 0.310 5.150 0.640 ;
        RECT  5.005 1.535 5.105 1.695 ;
        RECT  2.495 2.280 5.105 2.440 ;
        RECT  4.355 0.480 4.990 0.640 ;
        RECT  4.665 1.160 4.825 2.100 ;
        RECT  3.455 1.940 4.665 2.100 ;
        RECT  4.195 0.310 4.355 0.640 ;
        RECT  1.950 0.310 4.195 0.470 ;
        RECT  3.965 1.600 4.020 1.760 ;
        RECT  3.965 0.650 4.015 0.980 ;
        RECT  3.755 0.650 3.965 1.760 ;
        RECT  3.455 0.650 3.505 0.810 ;
        RECT  3.295 0.650 3.455 2.100 ;
        RECT  3.245 0.650 3.295 0.810 ;
        RECT  2.380 0.650 2.505 0.810 ;
        RECT  2.380 1.840 2.495 2.440 ;
        RECT  2.200 0.650 2.380 2.440 ;
        RECT  1.535 1.285 2.200 1.545 ;
        RECT  1.790 0.310 1.950 0.975 ;
        RECT  1.350 0.815 1.790 0.975 ;
        RECT  1.350 1.740 1.635 2.000 ;
        RECT  1.345 0.310 1.605 0.610 ;
        RECT  1.145 0.815 1.350 2.000 ;
        RECT  0.385 0.430 1.345 0.610 ;
        RECT  1.065 0.815 1.145 0.975 ;
        RECT  0.310 0.430 0.385 1.025 ;
        RECT  0.310 1.835 0.385 2.095 ;
        RECT  0.125 0.430 0.310 2.095 ;
    END
END DFFNSRHX8MTH

MACRO DFFQNX1MTH
    CLASS CORE ;
    FOREIGN DFFQNX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.115 0.720 7.280 2.120 ;
        RECT  6.995 0.720 7.115 0.980 ;
        RECT  7.025 1.685 7.115 2.120 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.700 2.615 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 -0.130 7.380 0.130 ;
        RECT  5.965 -0.130 6.565 0.250 ;
        RECT  4.565 -0.130 5.965 0.130 ;
        RECT  3.725 -0.130 4.565 0.325 ;
        RECT  1.065 -0.130 3.725 0.130 ;
        RECT  0.125 -0.130 1.065 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 2.740 7.380 3.000 ;
        RECT  6.060 2.570 6.660 3.000 ;
        RECT  4.480 2.740 6.060 3.000 ;
        RECT  4.220 2.620 4.480 3.000 ;
        RECT  3.620 2.740 4.220 3.000 ;
        RECT  3.020 2.620 3.620 3.000 ;
        RECT  2.200 2.740 3.020 3.000 ;
        RECT  1.940 2.620 2.200 3.000 ;
        RECT  0.555 2.740 1.940 3.000 ;
        RECT  0.295 2.205 0.555 3.000 ;
        RECT  0.000 2.740 0.295 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.845 1.215 6.935 1.475 ;
        RECT  6.685 1.215 6.845 2.115 ;
        RECT  6.250 1.955 6.685 2.115 ;
        RECT  6.345 0.430 6.505 1.390 ;
        RECT  5.695 0.430 6.345 0.590 ;
        RECT  6.295 1.130 6.345 1.390 ;
        RECT  6.035 1.930 6.250 2.115 ;
        RECT  6.035 0.790 6.135 0.950 ;
        RECT  5.875 0.790 6.035 2.115 ;
        RECT  5.830 1.510 5.875 1.770 ;
        RECT  5.555 0.430 5.695 1.300 ;
        RECT  5.535 0.430 5.555 2.475 ;
        RECT  4.865 0.430 5.535 0.590 ;
        RECT  5.395 1.140 5.535 2.475 ;
        RECT  5.100 2.315 5.395 2.475 ;
        RECT  5.215 0.800 5.355 0.960 ;
        RECT  5.055 0.800 5.215 2.105 ;
        RECT  4.980 1.845 5.055 2.105 ;
        RECT  4.915 1.945 4.980 2.105 ;
        RECT  4.755 1.945 4.915 2.440 ;
        RECT  4.715 1.360 4.875 1.620 ;
        RECT  4.045 2.280 4.755 2.440 ;
        RECT  4.190 1.360 4.715 1.520 ;
        RECT  4.315 1.915 4.575 2.100 ;
        RECT  3.615 1.940 4.315 2.100 ;
        RECT  3.930 1.360 4.190 1.760 ;
        RECT  3.785 2.280 4.045 2.540 ;
        RECT  3.840 1.360 3.930 1.520 ;
        RECT  3.680 0.680 3.840 1.520 ;
        RECT  2.770 2.280 3.785 2.440 ;
        RECT  3.540 0.680 3.680 0.840 ;
        RECT  3.455 1.805 3.615 2.100 ;
        RECT  3.380 0.310 3.540 0.840 ;
        RECT  3.200 1.805 3.455 1.965 ;
        RECT  1.280 0.310 3.380 0.470 ;
        RECT  3.040 0.805 3.200 1.965 ;
        RECT  1.830 1.355 3.040 1.515 ;
        RECT  2.880 1.805 3.040 1.965 ;
        RECT  2.670 0.670 2.830 1.165 ;
        RECT  2.495 2.280 2.770 2.475 ;
        RECT  1.385 1.005 2.670 1.165 ;
        RECT  1.635 2.280 2.495 2.440 ;
        RECT  0.970 0.665 2.490 0.825 ;
        RECT  1.375 2.280 1.635 2.515 ;
        RECT  1.385 1.935 1.435 2.095 ;
        RECT  1.225 1.005 1.385 2.095 ;
        RECT  0.995 2.280 1.375 2.440 ;
        RECT  0.910 1.005 1.225 1.165 ;
        RECT  1.175 1.935 1.225 2.095 ;
        RECT  0.835 1.375 0.995 2.440 ;
        RECT  0.730 0.525 0.970 0.825 ;
        RECT  0.730 1.375 0.835 1.535 ;
        RECT  0.710 0.525 0.730 1.535 ;
        RECT  0.570 0.665 0.710 1.535 ;
    END
END DFFQNX1MTH

MACRO DFFQNX2MTH
    CLASS CORE ;
    FOREIGN DFFQNX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.115 0.425 7.280 2.285 ;
        RECT  6.995 0.425 7.115 1.025 ;
        RECT  7.005 1.685 7.115 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.700 2.615 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 -0.130 7.380 0.130 ;
        RECT  5.965 -0.130 6.565 0.250 ;
        RECT  4.565 -0.130 5.965 0.130 ;
        RECT  3.725 -0.130 4.565 0.325 ;
        RECT  1.065 -0.130 3.725 0.130 ;
        RECT  0.125 -0.130 1.065 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 2.740 7.380 3.000 ;
        RECT  6.060 2.570 6.660 3.000 ;
        RECT  4.480 2.740 6.060 3.000 ;
        RECT  4.220 2.620 4.480 3.000 ;
        RECT  3.605 2.740 4.220 3.000 ;
        RECT  3.005 2.620 3.605 3.000 ;
        RECT  2.185 2.740 3.005 3.000 ;
        RECT  1.925 2.620 2.185 3.000 ;
        RECT  0.510 2.740 1.925 3.000 ;
        RECT  0.250 2.205 0.510 3.000 ;
        RECT  0.000 2.740 0.250 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.825 1.215 6.935 1.475 ;
        RECT  6.665 1.215 6.825 2.090 ;
        RECT  6.035 1.930 6.665 2.090 ;
        RECT  6.325 0.430 6.485 1.415 ;
        RECT  5.695 0.430 6.325 0.590 ;
        RECT  6.295 1.130 6.325 1.390 ;
        RECT  6.035 0.790 6.135 0.950 ;
        RECT  5.875 0.790 6.035 2.090 ;
        RECT  5.830 1.510 5.875 1.770 ;
        RECT  5.545 0.430 5.695 1.300 ;
        RECT  5.535 0.430 5.545 2.475 ;
        RECT  4.865 0.430 5.535 0.590 ;
        RECT  5.385 1.140 5.535 2.475 ;
        RECT  5.100 2.315 5.385 2.475 ;
        RECT  5.205 0.800 5.355 0.960 ;
        RECT  5.045 0.800 5.205 2.105 ;
        RECT  4.980 1.845 5.045 2.105 ;
        RECT  4.915 1.945 4.980 2.105 ;
        RECT  4.755 1.945 4.915 2.440 ;
        RECT  4.705 1.360 4.865 1.620 ;
        RECT  4.045 2.280 4.755 2.440 ;
        RECT  4.180 1.360 4.705 1.520 ;
        RECT  4.315 1.915 4.575 2.100 ;
        RECT  3.615 1.940 4.315 2.100 ;
        RECT  3.920 1.360 4.180 1.760 ;
        RECT  3.785 2.280 4.045 2.540 ;
        RECT  3.840 1.360 3.920 1.520 ;
        RECT  3.680 0.680 3.840 1.520 ;
        RECT  2.755 2.280 3.785 2.440 ;
        RECT  3.540 0.680 3.680 0.840 ;
        RECT  3.455 1.805 3.615 2.100 ;
        RECT  3.380 0.310 3.540 0.840 ;
        RECT  3.200 1.805 3.455 1.965 ;
        RECT  1.280 0.310 3.380 0.470 ;
        RECT  3.040 0.805 3.200 1.965 ;
        RECT  1.815 1.355 3.040 1.515 ;
        RECT  2.865 1.805 3.040 1.965 ;
        RECT  2.670 0.670 2.830 1.165 ;
        RECT  2.495 2.280 2.755 2.475 ;
        RECT  1.340 1.005 2.670 1.165 ;
        RECT  1.590 2.280 2.495 2.440 ;
        RECT  0.970 0.665 2.490 0.825 ;
        RECT  1.330 2.280 1.590 2.515 ;
        RECT  1.340 1.935 1.390 2.095 ;
        RECT  1.180 1.005 1.340 2.095 ;
        RECT  0.950 2.280 1.330 2.440 ;
        RECT  0.910 1.005 1.180 1.165 ;
        RECT  1.130 1.935 1.180 2.095 ;
        RECT  0.730 0.525 0.970 0.825 ;
        RECT  0.790 1.375 0.950 2.440 ;
        RECT  0.730 1.375 0.790 1.535 ;
        RECT  0.710 0.525 0.730 1.535 ;
        RECT  0.570 0.665 0.710 1.535 ;
    END
END DFFQNX2MTH

MACRO DFFQNX4MTH
    CLASS CORE ;
    FOREIGN DFFQNX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.280 0.425 7.315 2.015 ;
        RECT  7.135 0.425 7.280 2.285 ;
        RECT  6.995 0.425 7.135 1.025 ;
        RECT  7.005 1.685 7.135 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.700 2.615 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 -0.130 7.790 0.130 ;
        RECT  5.965 -0.130 6.565 0.250 ;
        RECT  4.565 -0.130 5.965 0.130 ;
        RECT  3.725 -0.130 4.565 0.325 ;
        RECT  1.065 -0.130 3.725 0.130 ;
        RECT  0.125 -0.130 1.065 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 2.740 7.790 3.000 ;
        RECT  6.060 2.570 6.660 3.000 ;
        RECT  4.480 2.740 6.060 3.000 ;
        RECT  4.220 2.620 4.480 3.000 ;
        RECT  3.605 2.740 4.220 3.000 ;
        RECT  3.005 2.620 3.605 3.000 ;
        RECT  2.185 2.740 3.005 3.000 ;
        RECT  1.925 2.620 2.185 3.000 ;
        RECT  0.515 2.740 1.925 3.000 ;
        RECT  0.255 2.205 0.515 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.825 1.215 6.955 1.475 ;
        RECT  6.665 1.215 6.825 2.105 ;
        RECT  6.035 1.945 6.665 2.105 ;
        RECT  6.315 0.430 6.475 1.405 ;
        RECT  5.695 0.430 6.315 0.590 ;
        RECT  6.035 0.815 6.135 0.975 ;
        RECT  5.875 0.815 6.035 2.105 ;
        RECT  5.780 1.525 5.875 1.785 ;
        RECT  5.535 0.430 5.695 1.300 ;
        RECT  4.865 0.430 5.535 0.590 ;
        RECT  5.490 1.140 5.535 1.300 ;
        RECT  5.330 1.140 5.490 2.465 ;
        RECT  5.150 0.800 5.355 0.960 ;
        RECT  5.100 2.305 5.330 2.465 ;
        RECT  4.990 0.800 5.150 2.105 ;
        RECT  4.950 1.845 4.990 2.105 ;
        RECT  4.915 1.945 4.950 2.105 ;
        RECT  4.755 1.945 4.915 2.440 ;
        RECT  4.650 1.360 4.810 1.620 ;
        RECT  4.045 2.280 4.755 2.440 ;
        RECT  4.180 1.360 4.650 1.520 ;
        RECT  4.315 1.915 4.575 2.100 ;
        RECT  3.615 1.940 4.315 2.100 ;
        RECT  3.920 1.360 4.180 1.760 ;
        RECT  3.785 2.280 4.045 2.540 ;
        RECT  3.840 1.360 3.920 1.520 ;
        RECT  3.680 0.680 3.840 1.520 ;
        RECT  2.755 2.280 3.785 2.440 ;
        RECT  3.540 0.680 3.680 0.840 ;
        RECT  3.455 1.805 3.615 2.100 ;
        RECT  3.380 0.310 3.540 0.840 ;
        RECT  3.200 1.805 3.455 1.965 ;
        RECT  1.280 0.310 3.380 0.470 ;
        RECT  3.040 0.805 3.200 1.965 ;
        RECT  1.815 1.355 3.040 1.515 ;
        RECT  2.865 1.805 3.040 1.965 ;
        RECT  2.670 0.670 2.830 1.165 ;
        RECT  2.495 2.280 2.755 2.475 ;
        RECT  1.345 1.005 2.670 1.165 ;
        RECT  1.745 2.280 2.495 2.440 ;
        RECT  0.970 0.665 2.490 0.825 ;
        RECT  1.585 2.280 1.745 2.485 ;
        RECT  0.955 2.325 1.585 2.485 ;
        RECT  1.345 1.955 1.395 2.115 ;
        RECT  1.185 1.005 1.345 2.115 ;
        RECT  0.910 1.005 1.185 1.165 ;
        RECT  1.135 1.955 1.185 2.115 ;
        RECT  0.730 0.525 0.970 0.825 ;
        RECT  0.795 1.375 0.955 2.485 ;
        RECT  0.730 1.375 0.795 1.535 ;
        RECT  0.710 0.525 0.730 1.535 ;
        RECT  0.570 0.665 0.710 1.535 ;
    END
END DFFQNX4MTH

MACRO DFFQX1MTH
    CLASS CORE ;
    FOREIGN DFFQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.250 1.290 7.280 1.580 ;
        RECT  6.990 0.735 7.250 2.015 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.700 2.565 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.960 -0.130 7.380 0.130 ;
        RECT  6.020 -0.130 6.960 0.250 ;
        RECT  4.710 -0.130 6.020 0.130 ;
        RECT  4.370 -0.130 4.710 0.325 ;
        RECT  4.110 -0.130 4.370 0.665 ;
        RECT  3.770 -0.130 4.110 0.325 ;
        RECT  0.395 -0.130 3.770 0.130 ;
        RECT  0.135 -0.130 0.395 0.325 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.970 2.740 7.380 3.000 ;
        RECT  6.030 2.555 6.970 3.000 ;
        RECT  4.540 2.740 6.030 3.000 ;
        RECT  4.280 2.620 4.540 3.000 ;
        RECT  3.645 2.740 4.280 3.000 ;
        RECT  3.045 2.620 3.645 3.000 ;
        RECT  2.135 2.740 3.045 3.000 ;
        RECT  1.875 2.620 2.135 3.000 ;
        RECT  0.385 2.740 1.875 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.650 1.230 6.770 1.490 ;
        RECT  6.490 0.445 6.650 2.305 ;
        RECT  5.260 0.445 6.490 0.605 ;
        RECT  5.340 2.145 6.490 2.305 ;
        RECT  6.075 0.815 6.280 1.025 ;
        RECT  6.075 1.685 6.280 1.945 ;
        RECT  5.915 0.815 6.075 1.945 ;
        RECT  5.815 1.210 5.915 1.470 ;
        RECT  5.540 0.820 5.590 1.080 ;
        RECT  5.380 0.820 5.540 1.865 ;
        RECT  5.330 0.820 5.380 1.080 ;
        RECT  5.000 1.705 5.380 1.865 ;
        RECT  5.180 2.045 5.340 2.305 ;
        RECT  5.000 0.445 5.260 0.640 ;
        RECT  4.170 1.220 5.050 1.380 ;
        RECT  4.840 1.705 5.000 2.440 ;
        RECT  4.085 2.280 4.840 2.440 ;
        RECT  4.400 1.675 4.660 2.100 ;
        RECT  3.615 1.940 4.400 2.100 ;
        RECT  3.910 1.220 4.170 1.760 ;
        RECT  3.825 2.280 4.085 2.535 ;
        RECT  3.750 1.220 3.910 1.380 ;
        RECT  2.755 2.280 3.825 2.440 ;
        RECT  3.590 0.630 3.750 1.380 ;
        RECT  3.455 1.805 3.615 2.100 ;
        RECT  3.430 0.325 3.590 0.890 ;
        RECT  3.200 1.805 3.455 1.965 ;
        RECT  1.280 0.325 3.430 0.485 ;
        RECT  3.040 0.805 3.200 1.965 ;
        RECT  1.700 1.355 3.040 1.515 ;
        RECT  2.815 1.805 3.040 1.965 ;
        RECT  2.670 0.670 2.830 1.165 ;
        RECT  2.445 2.280 2.755 2.475 ;
        RECT  1.255 1.005 2.670 1.165 ;
        RECT  0.940 0.665 2.490 0.825 ;
        RECT  1.615 2.280 2.445 2.440 ;
        RECT  1.455 2.280 1.615 2.485 ;
        RECT  0.730 2.325 1.455 2.485 ;
        RECT  1.255 1.940 1.305 2.100 ;
        RECT  1.095 1.005 1.255 2.100 ;
        RECT  0.910 1.005 1.095 1.165 ;
        RECT  1.045 1.940 1.095 2.100 ;
        RECT  0.730 0.415 0.940 0.825 ;
        RECT  0.680 0.415 0.730 2.485 ;
        RECT  0.570 0.665 0.680 2.485 ;
    END
END DFFQX1MTH

MACRO DFFQX2MTH
    CLASS CORE ;
    FOREIGN DFFQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.250 1.290 7.280 1.580 ;
        RECT  6.990 0.425 7.250 2.300 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.700 2.565 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.710 -0.130 7.380 0.130 ;
        RECT  6.110 -0.130 6.710 0.250 ;
        RECT  4.370 -0.130 6.110 0.130 ;
        RECT  4.110 -0.130 4.370 0.665 ;
        RECT  3.770 -0.130 4.110 0.325 ;
        RECT  0.395 -0.130 3.770 0.130 ;
        RECT  0.135 -0.130 0.395 0.325 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.630 2.740 7.380 3.000 ;
        RECT  6.030 2.575 6.630 3.000 ;
        RECT  4.540 2.740 6.030 3.000 ;
        RECT  4.280 2.620 4.540 3.000 ;
        RECT  3.600 2.740 4.280 3.000 ;
        RECT  3.000 2.620 3.600 3.000 ;
        RECT  2.135 2.740 3.000 3.000 ;
        RECT  1.875 2.620 2.135 3.000 ;
        RECT  0.385 2.740 1.875 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.650 1.230 6.770 1.490 ;
        RECT  6.490 0.455 6.650 2.325 ;
        RECT  5.000 0.455 6.490 0.615 ;
        RECT  5.340 2.165 6.490 2.325 ;
        RECT  6.075 0.815 6.280 0.975 ;
        RECT  6.075 1.685 6.280 1.945 ;
        RECT  5.915 0.815 6.075 1.945 ;
        RECT  5.815 1.210 5.915 1.470 ;
        RECT  5.540 0.820 5.590 1.080 ;
        RECT  5.380 0.820 5.540 1.825 ;
        RECT  5.330 0.820 5.380 1.080 ;
        RECT  5.000 1.665 5.380 1.825 ;
        RECT  5.180 2.165 5.340 2.425 ;
        RECT  4.790 1.180 5.050 1.410 ;
        RECT  4.840 1.665 5.000 2.440 ;
        RECT  4.085 2.280 4.840 2.440 ;
        RECT  4.170 1.250 4.790 1.410 ;
        RECT  4.400 1.685 4.660 2.100 ;
        RECT  3.615 1.940 4.400 2.100 ;
        RECT  3.910 1.250 4.170 1.760 ;
        RECT  3.825 2.280 4.085 2.540 ;
        RECT  3.750 1.250 3.910 1.410 ;
        RECT  2.755 2.280 3.825 2.440 ;
        RECT  3.590 0.630 3.750 1.410 ;
        RECT  3.455 1.805 3.615 2.100 ;
        RECT  3.430 0.325 3.590 0.890 ;
        RECT  3.200 1.805 3.455 1.965 ;
        RECT  1.280 0.325 3.430 0.485 ;
        RECT  3.040 0.805 3.200 1.965 ;
        RECT  1.725 1.355 3.040 1.515 ;
        RECT  2.815 1.805 3.040 1.965 ;
        RECT  2.670 0.670 2.830 1.165 ;
        RECT  2.445 2.280 2.755 2.475 ;
        RECT  1.255 1.005 2.670 1.165 ;
        RECT  0.940 0.665 2.490 0.825 ;
        RECT  1.615 2.280 2.445 2.440 ;
        RECT  1.455 2.280 1.615 2.465 ;
        RECT  0.730 2.305 1.455 2.465 ;
        RECT  1.255 1.925 1.305 2.085 ;
        RECT  1.095 1.005 1.255 2.085 ;
        RECT  0.910 1.005 1.095 1.165 ;
        RECT  1.045 1.925 1.095 2.085 ;
        RECT  0.730 0.415 0.940 0.825 ;
        RECT  0.680 0.415 0.730 2.465 ;
        RECT  0.570 0.665 0.680 2.465 ;
    END
END DFFQX2MTH

MACRO DFFQX4MTH
    CLASS CORE ;
    FOREIGN DFFQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.040 0.425 7.300 2.300 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 1.670 2.720 1.975 ;
        END
        AntennaGateArea 0.104 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.710 -0.130 7.790 0.130 ;
        RECT  6.110 -0.130 6.710 0.250 ;
        RECT  4.370 -0.130 6.110 0.130 ;
        RECT  4.110 -0.130 4.370 0.665 ;
        RECT  3.770 -0.130 4.110 0.325 ;
        RECT  0.395 -0.130 3.770 0.130 ;
        RECT  0.135 -0.130 0.395 0.325 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.630 2.740 7.790 3.000 ;
        RECT  6.030 2.575 6.630 3.000 ;
        RECT  4.540 2.740 6.030 3.000 ;
        RECT  4.280 2.620 4.540 3.000 ;
        RECT  3.595 2.740 4.280 3.000 ;
        RECT  2.995 2.620 3.595 3.000 ;
        RECT  1.920 2.740 2.995 3.000 ;
        RECT  1.660 2.620 1.920 3.000 ;
        RECT  0.385 2.740 1.660 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.650 1.230 6.860 1.490 ;
        RECT  6.490 0.465 6.650 2.395 ;
        RECT  5.000 0.465 6.490 0.625 ;
        RECT  6.360 1.230 6.490 1.490 ;
        RECT  5.340 2.235 6.490 2.395 ;
        RECT  6.075 0.815 6.280 0.975 ;
        RECT  6.075 1.685 6.280 1.945 ;
        RECT  5.915 0.815 6.075 1.945 ;
        RECT  5.815 1.210 5.915 1.470 ;
        RECT  5.540 0.805 5.590 1.065 ;
        RECT  5.380 0.805 5.540 1.785 ;
        RECT  5.330 0.805 5.380 1.065 ;
        RECT  5.000 1.625 5.380 1.785 ;
        RECT  5.180 2.235 5.340 2.495 ;
        RECT  4.170 1.145 5.050 1.305 ;
        RECT  4.840 1.625 5.000 2.440 ;
        RECT  4.085 2.280 4.840 2.440 ;
        RECT  4.400 1.575 4.660 2.100 ;
        RECT  3.615 1.940 4.400 2.100 ;
        RECT  3.910 1.145 4.170 1.760 ;
        RECT  3.825 2.280 4.085 2.535 ;
        RECT  3.750 1.145 3.910 1.305 ;
        RECT  2.460 2.280 3.825 2.440 ;
        RECT  3.590 0.575 3.750 1.305 ;
        RECT  3.455 1.805 3.615 2.100 ;
        RECT  3.430 0.310 3.590 0.835 ;
        RECT  3.200 1.805 3.455 1.965 ;
        RECT  1.280 0.310 3.430 0.470 ;
        RECT  3.040 0.825 3.200 1.965 ;
        RECT  1.590 1.330 3.040 1.490 ;
        RECT  2.905 1.805 3.040 1.965 ;
        RECT  2.670 0.670 2.830 1.150 ;
        RECT  1.070 0.990 2.670 1.150 ;
        RECT  0.940 0.650 2.490 0.810 ;
        RECT  2.200 2.180 2.460 2.440 ;
        RECT  1.445 2.280 2.200 2.440 ;
        RECT  1.285 2.280 1.445 2.470 ;
        RECT  0.730 2.310 1.285 2.470 ;
        RECT  1.070 1.860 1.120 2.120 ;
        RECT  0.910 0.990 1.070 2.120 ;
        RECT  0.730 0.510 0.940 0.810 ;
        RECT  0.680 0.510 0.730 2.470 ;
        RECT  0.570 0.650 0.680 2.470 ;
    END
END DFFQX4MTH

MACRO DFFRHQX1MTH
    CLASS CORE ;
    FOREIGN DFFRHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.285 5.400 1.730 ;
        END
        AntennaGateArea 0.143 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.045 1.370 10.150 2.045 ;
        RECT  10.045 0.735 10.075 0.995 ;
        RECT  9.885 0.735 10.045 2.045 ;
        END
        AntennaDiffArea 0.362 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.470 1.030 2.770 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.475 1.145 0.800 1.580 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.020 -0.130 10.250 0.130 ;
        RECT  9.860 -0.130 10.020 0.300 ;
        RECT  9.555 -0.130 9.860 0.130 ;
        RECT  8.955 -0.130 9.555 0.425 ;
        RECT  8.735 -0.130 8.955 0.130 ;
        RECT  8.135 -0.130 8.735 0.425 ;
        RECT  5.245 -0.130 8.135 0.130 ;
        RECT  4.985 -0.130 5.245 0.415 ;
        RECT  2.125 -0.130 4.985 0.130 ;
        RECT  1.965 -0.130 2.125 0.300 ;
        RECT  0.605 -0.130 1.965 0.130 ;
        RECT  0.330 -0.130 0.605 0.345 ;
        RECT  0.000 -0.130 0.330 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.520 2.740 10.250 3.000 ;
        RECT  8.880 2.425 9.520 3.000 ;
        RECT  7.630 2.740 8.880 3.000 ;
        RECT  7.370 2.520 7.630 3.000 ;
        RECT  1.945 2.740 7.370 3.000 ;
        RECT  1.685 2.570 1.945 3.000 ;
        RECT  0.790 2.740 1.685 3.000 ;
        RECT  0.265 2.230 0.790 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.440 1.215 9.705 1.475 ;
        RECT  9.280 1.215 9.440 2.240 ;
        RECT  9.205 1.215 9.280 1.475 ;
        RECT  8.210 2.080 9.280 2.240 ;
        RECT  8.805 1.735 9.100 1.895 ;
        RECT  8.805 0.765 9.035 1.025 ;
        RECT  8.775 0.765 8.805 1.895 ;
        RECT  8.645 0.855 8.775 1.895 ;
        RECT  8.520 1.160 8.645 1.760 ;
        RECT  8.120 1.505 8.250 1.765 ;
        RECT  7.950 2.080 8.210 2.515 ;
        RECT  7.990 0.605 8.120 1.765 ;
        RECT  7.960 0.605 7.990 1.600 ;
        RECT  7.955 0.605 7.960 0.765 ;
        RECT  7.795 0.310 7.955 0.765 ;
        RECT  7.615 2.080 7.950 2.240 ;
        RECT  6.560 0.310 7.795 0.470 ;
        RECT  7.455 0.785 7.615 2.240 ;
        RECT  6.900 0.785 7.455 0.945 ;
        RECT  7.190 1.815 7.455 2.075 ;
        RECT  7.010 1.475 7.225 1.635 ;
        RECT  6.850 1.475 7.010 2.560 ;
        RECT  6.740 0.665 6.900 0.945 ;
        RECT  3.885 2.400 6.850 2.560 ;
        RECT  6.560 1.145 6.745 1.305 ;
        RECT  6.220 1.960 6.670 2.220 ;
        RECT  6.400 0.310 6.560 1.305 ;
        RECT  5.740 0.310 6.400 0.470 ;
        RECT  6.060 0.665 6.220 2.220 ;
        RECT  5.950 0.665 6.060 0.925 ;
        RECT  4.840 2.060 6.060 2.220 ;
        RECT  5.740 1.330 5.880 1.590 ;
        RECT  5.580 0.310 5.740 0.755 ;
        RECT  5.580 0.940 5.740 1.590 ;
        RECT  4.735 0.595 5.580 0.755 ;
        RECT  4.395 0.940 5.580 1.100 ;
        RECT  4.680 1.385 4.840 2.220 ;
        RECT  4.575 0.310 4.735 0.755 ;
        RECT  2.465 0.310 4.575 0.470 ;
        RECT  4.235 0.725 4.395 2.170 ;
        RECT  4.065 2.010 4.235 2.170 ;
        RECT  3.885 1.050 3.985 1.210 ;
        RECT  3.725 0.680 3.885 1.210 ;
        RECT  3.725 1.425 3.885 2.560 ;
        RECT  3.110 0.680 3.725 0.840 ;
        RECT  3.545 1.425 3.725 1.585 ;
        RECT  2.285 2.400 3.725 2.560 ;
        RECT  3.385 1.125 3.545 1.585 ;
        RECT  3.385 1.765 3.545 2.220 ;
        RECT  3.295 1.125 3.385 1.385 ;
        RECT  2.625 2.060 3.385 2.220 ;
        RECT  2.950 0.680 3.110 1.810 ;
        RECT  2.655 0.680 2.950 0.840 ;
        RECT  2.465 1.760 2.625 2.220 ;
        RECT  2.305 0.310 2.465 0.840 ;
        RECT  2.015 1.760 2.465 1.920 ;
        RECT  1.845 0.680 2.305 0.840 ;
        RECT  2.125 2.230 2.285 2.560 ;
        RECT  1.665 2.230 2.125 2.390 ;
        RECT  1.845 1.550 2.015 1.920 ;
        RECT  1.685 0.680 1.845 1.920 ;
        RECT  1.505 0.310 1.765 0.495 ;
        RECT  1.635 0.680 1.685 0.840 ;
        RECT  1.320 1.550 1.685 1.810 ;
        RECT  1.405 2.110 1.665 2.390 ;
        RECT  0.945 0.335 1.505 0.495 ;
        RECT  1.140 2.230 1.405 2.390 ;
        RECT  1.140 0.680 1.385 1.025 ;
        RECT  1.125 0.680 1.140 2.390 ;
        RECT  0.980 0.865 1.125 2.390 ;
        RECT  0.785 0.335 0.945 0.685 ;
        RECT  0.335 0.525 0.785 0.685 ;
        RECT  0.285 1.770 0.385 1.930 ;
        RECT  0.285 0.525 0.335 0.890 ;
        RECT  0.125 0.525 0.285 1.930 ;
    END
END DFFRHQX1MTH

MACRO DFFRHQX2MTH
    CLASS CORE ;
    FOREIGN DFFRHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.785 1.330 7.780 1.490 ;
        RECT  6.645 1.330 6.785 1.540 ;
        RECT  6.485 1.330 6.645 1.710 ;
        RECT  5.855 1.550 6.485 1.710 ;
        RECT  5.640 1.550 5.855 1.795 ;
        RECT  5.595 1.290 5.640 1.795 ;
        RECT  5.430 1.290 5.595 1.710 ;
        END
        AntennaGateArea 0.1781 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.710 0.745 10.915 2.375 ;
        RECT  10.360 0.745 10.710 0.905 ;
        RECT  10.580 1.700 10.710 2.375 ;
        RECT  10.350 1.700 10.580 1.990 ;
        RECT  10.200 0.380 10.360 0.905 ;
        END
        AntennaDiffArea 0.426 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.415 1.005 2.575 1.255 ;
        RECT  2.150 0.880 2.415 1.255 ;
        RECT  2.070 1.005 2.150 1.255 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.135 0.785 1.580 ;
        END
        AntennaGateArea 0.143 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.920 -0.130 11.070 0.130 ;
        RECT  10.660 -0.130 10.920 0.565 ;
        RECT  9.810 -0.130 10.660 0.130 ;
        RECT  9.650 -0.130 9.810 0.520 ;
        RECT  5.445 -0.130 9.650 0.130 ;
        RECT  4.845 -0.130 5.445 0.405 ;
        RECT  0.950 -0.130 4.845 0.130 ;
        RECT  0.485 -0.130 0.950 0.250 ;
        RECT  0.325 -0.130 0.485 0.480 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.220 2.740 11.070 3.000 ;
        RECT  9.775 2.555 10.220 3.000 ;
        RECT  8.530 2.740 9.775 3.000 ;
        RECT  8.270 2.620 8.530 3.000 ;
        RECT  3.830 2.740 8.270 3.000 ;
        RECT  3.670 2.570 3.830 3.000 ;
        RECT  0.815 2.740 3.670 3.000 ;
        RECT  0.215 2.280 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.160 1.150 10.530 1.410 ;
        RECT  10.000 1.150 10.160 2.375 ;
        RECT  9.110 2.215 10.000 2.375 ;
        RECT  9.570 1.405 9.820 1.665 ;
        RECT  9.410 0.945 9.570 1.665 ;
        RECT  9.220 0.945 9.410 1.205 ;
        RECT  9.060 0.310 9.220 1.205 ;
        RECT  8.880 1.505 9.150 1.765 ;
        RECT  8.850 2.215 9.110 2.505 ;
        RECT  8.720 0.310 8.880 1.765 ;
        RECT  8.470 2.215 8.850 2.375 ;
        RECT  6.010 0.310 8.720 0.470 ;
        RECT  8.310 0.650 8.470 2.375 ;
        RECT  6.755 0.650 8.310 0.810 ;
        RECT  7.635 2.215 8.310 2.375 ;
        RECT  7.970 0.990 8.130 2.035 ;
        RECT  6.455 0.990 7.970 1.150 ;
        RECT  7.955 1.670 7.970 2.035 ;
        RECT  7.185 1.670 7.955 1.830 ;
        RECT  7.475 2.025 7.635 2.375 ;
        RECT  7.365 2.025 7.475 2.185 ;
        RECT  4.175 2.400 7.295 2.560 ;
        RECT  7.025 1.670 7.185 2.220 ;
        RECT  6.870 1.895 7.025 2.220 ;
        RECT  5.220 2.050 6.870 2.220 ;
        RECT  6.295 0.650 6.455 1.150 ;
        RECT  5.955 0.940 6.115 1.365 ;
        RECT  5.850 0.310 6.010 0.760 ;
        RECT  4.865 0.940 5.955 1.100 ;
        RECT  4.550 0.600 5.850 0.760 ;
        RECT  5.060 1.295 5.220 2.220 ;
        RECT  4.705 0.940 4.865 2.165 ;
        RECT  4.210 0.940 4.705 1.100 ;
        RECT  4.555 2.005 4.705 2.165 ;
        RECT  4.390 0.310 4.550 0.760 ;
        RECT  4.365 1.315 4.525 1.790 ;
        RECT  1.845 0.310 4.390 0.470 ;
        RECT  3.870 1.315 4.365 1.475 ;
        RECT  4.050 0.665 4.210 1.100 ;
        RECT  4.015 2.230 4.175 2.560 ;
        RECT  3.460 2.230 4.015 2.390 ;
        RECT  3.710 0.650 3.870 1.475 ;
        RECT  2.915 0.650 3.710 0.810 ;
        RECT  3.525 1.315 3.710 1.475 ;
        RECT  3.300 1.655 3.460 2.495 ;
        RECT  3.255 1.655 3.300 1.815 ;
        RECT  1.695 2.335 3.300 2.495 ;
        RECT  3.095 0.990 3.255 1.815 ;
        RECT  2.915 1.995 3.120 2.155 ;
        RECT  2.755 0.650 2.915 2.155 ;
        RECT  2.635 0.650 2.755 0.810 ;
        RECT  1.900 1.440 2.190 1.945 ;
        RECT  1.845 1.440 1.900 1.690 ;
        RECT  1.685 0.310 1.845 1.690 ;
        RECT  1.415 1.870 1.695 2.495 ;
        RECT  1.305 1.430 1.685 1.690 ;
        RECT  1.235 0.425 1.495 0.635 ;
        RECT  1.125 1.870 1.415 2.030 ;
        RECT  1.125 0.815 1.395 1.250 ;
        RECT  0.830 0.475 1.235 0.635 ;
        RECT  1.115 0.815 1.125 2.030 ;
        RECT  0.965 1.090 1.115 2.030 ;
        RECT  0.670 0.475 0.830 0.910 ;
        RECT  0.385 0.750 0.670 0.910 ;
        RECT  0.285 0.750 0.385 0.940 ;
        RECT  0.285 1.770 0.385 1.930 ;
        RECT  0.125 0.750 0.285 1.930 ;
    END
END DFFRHQX2MTH

MACRO DFFRHQX4MTH
    CLASS CORE ;
    FOREIGN DFFRHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.660 1.085 8.920 1.635 ;
        RECT  8.620 1.375 8.660 1.635 ;
        END
        AntennaGateArea 0.1703 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 0.385 10.970 2.405 ;
        RECT  10.660 0.385 10.730 0.985 ;
        RECT  10.660 1.805 10.730 2.405 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.880 2.900 1.380 ;
        END
        AntennaGateArea 0.1664 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.120 0.760 1.680 ;
        END
        AntennaGateArea 0.1612 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.330 -0.130 11.480 0.130 ;
        RECT  10.070 -0.130 10.330 0.515 ;
        RECT  9.715 -0.130 10.070 0.130 ;
        RECT  9.115 -0.130 9.715 0.515 ;
        RECT  6.085 -0.130 9.115 0.130 ;
        RECT  5.485 -0.130 6.085 0.460 ;
        RECT  2.680 -0.130 5.485 0.130 ;
        RECT  2.480 -0.130 2.680 0.680 ;
        RECT  0.680 -0.130 2.480 0.130 ;
        RECT  0.420 -0.130 0.680 0.300 ;
        RECT  0.000 -0.130 0.420 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.285 2.740 11.480 3.000 ;
        RECT  9.785 2.415 10.285 3.000 ;
        RECT  8.470 2.740 9.785 3.000 ;
        RECT  8.210 2.295 8.470 3.000 ;
        RECT  6.495 2.740 8.210 3.000 ;
        RECT  6.235 2.620 6.495 3.000 ;
        RECT  5.395 2.740 6.235 3.000 ;
        RECT  5.135 2.620 5.395 3.000 ;
        RECT  2.110 2.740 5.135 3.000 ;
        RECT  1.610 2.570 2.110 3.000 ;
        RECT  0.845 2.740 1.610 3.000 ;
        RECT  0.245 2.365 0.845 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.285 1.230 10.525 1.490 ;
        RECT  10.125 1.230 10.285 2.235 ;
        RECT  10.025 1.230 10.125 1.490 ;
        RECT  9.605 2.075 10.125 2.235 ;
        RECT  9.790 1.735 9.900 1.895 ;
        RECT  9.790 0.765 9.850 1.025 ;
        RECT  9.630 0.765 9.790 1.895 ;
        RECT  9.440 1.135 9.630 1.395 ;
        RECT  9.445 2.075 9.605 2.455 ;
        RECT  8.820 2.295 9.445 2.455 ;
        RECT  9.100 0.745 9.260 2.115 ;
        RECT  8.830 0.745 9.100 0.905 ;
        RECT  9.000 1.855 9.100 2.115 ;
        RECT  8.670 0.310 8.830 0.905 ;
        RECT  8.660 1.955 8.820 2.455 ;
        RECT  7.615 0.310 8.670 0.470 ;
        RECT  8.440 1.955 8.660 2.115 ;
        RECT  8.280 0.650 8.440 2.115 ;
        RECT  7.795 0.650 8.280 0.810 ;
        RECT  7.610 1.955 8.280 2.115 ;
        RECT  7.840 1.470 8.100 1.775 ;
        RECT  7.275 1.470 7.840 1.630 ;
        RECT  7.455 0.310 7.615 1.145 ;
        RECT  7.450 1.815 7.610 2.115 ;
        RECT  6.740 0.310 7.455 0.470 ;
        RECT  7.300 1.815 7.450 1.975 ;
        RECT  7.020 2.185 7.280 2.440 ;
        RECT  7.120 0.650 7.275 1.630 ;
        RECT  7.115 0.650 7.120 1.980 ;
        RECT  7.015 0.650 7.115 0.810 ;
        RECT  6.960 1.470 7.115 1.980 ;
        RECT  4.955 2.280 7.020 2.440 ;
        RECT  6.840 1.720 6.960 1.980 ;
        RECT  6.695 0.990 6.855 1.315 ;
        RECT  6.680 1.720 6.840 2.100 ;
        RECT  6.580 0.310 6.740 0.810 ;
        RECT  6.115 0.990 6.695 1.150 ;
        RECT  5.245 1.940 6.680 2.100 ;
        RECT  4.920 0.650 6.580 0.810 ;
        RECT  5.515 0.990 6.115 1.760 ;
        RECT  4.605 0.990 5.515 1.150 ;
        RECT  5.085 1.455 5.245 2.100 ;
        RECT  4.795 2.280 4.955 2.560 ;
        RECT  4.760 0.365 4.920 0.810 ;
        RECT  4.255 2.400 4.795 2.560 ;
        RECT  3.580 0.650 4.760 0.810 ;
        RECT  4.445 0.990 4.605 2.210 ;
        RECT  3.240 0.310 4.455 0.470 ;
        RECT  4.095 1.165 4.255 2.560 ;
        RECT  3.920 1.165 4.095 1.325 ;
        RECT  2.495 2.400 4.095 2.560 ;
        RECT  3.760 1.065 3.920 1.325 ;
        RECT  3.580 1.545 3.895 1.805 ;
        RECT  3.420 0.650 3.580 2.220 ;
        RECT  2.865 2.060 3.420 2.220 ;
        RECT  3.080 0.310 3.240 1.880 ;
        RECT  3.050 0.435 3.080 0.695 ;
        RECT  3.050 1.620 3.080 1.880 ;
        RECT  2.705 1.600 2.865 2.220 ;
        RECT  2.155 1.600 2.705 1.760 ;
        RECT  2.335 2.055 2.495 2.560 ;
        RECT  1.790 2.055 2.335 2.215 ;
        RECT  1.020 0.310 2.300 0.470 ;
        RECT  1.995 0.680 2.155 1.760 ;
        RECT  1.760 0.680 1.995 0.840 ;
        RECT  1.570 1.600 1.995 1.760 ;
        RECT  1.530 2.055 1.790 2.270 ;
        RECT  1.410 1.470 1.570 1.760 ;
        RECT  1.105 2.055 1.530 2.215 ;
        RECT  1.410 0.680 1.510 0.840 ;
        RECT  1.250 0.680 1.410 1.280 ;
        RECT  1.105 1.120 1.250 1.280 ;
        RECT  0.945 1.120 1.105 2.215 ;
        RECT  0.860 0.310 1.020 0.925 ;
        RECT  0.355 0.765 0.860 0.925 ;
        RECT  0.330 1.790 0.360 2.050 ;
        RECT  0.330 0.765 0.355 1.025 ;
        RECT  0.170 0.765 0.330 2.050 ;
    END
END DFFRHQX4MTH

MACRO DFFRHQX8MTH
    CLASS CORE ;
    FOREIGN DFFRHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.660 1.085 8.920 1.635 ;
        RECT  8.620 1.375 8.660 1.635 ;
        END
        AntennaGateArea 0.1703 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 0.385 11.705 2.405 ;
        RECT  10.950 1.085 11.355 1.785 ;
        RECT  10.600 0.385 10.950 2.405 ;
        RECT  10.470 0.385 10.600 0.985 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.285 0.880 2.835 1.380 ;
        END
        AntennaGateArea 0.1664 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.120 0.760 1.695 ;
        END
        AntennaGateArea 0.1612 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 -0.130 12.300 0.130 ;
        RECT  11.915 -0.130 12.175 0.985 ;
        RECT  10.185 -0.130 11.915 0.130 ;
        RECT  9.925 -0.130 10.185 0.515 ;
        RECT  9.670 -0.130 9.925 0.130 ;
        RECT  9.070 -0.130 9.670 0.515 ;
        RECT  6.085 -0.130 9.070 0.130 ;
        RECT  5.485 -0.130 6.085 0.460 ;
        RECT  2.590 -0.130 5.485 0.130 ;
        RECT  2.330 -0.130 2.590 0.680 ;
        RECT  0.680 -0.130 2.330 0.130 ;
        RECT  0.420 -0.130 0.680 0.300 ;
        RECT  0.000 -0.130 0.420 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.200 2.740 12.300 3.000 ;
        RECT  9.780 2.415 10.200 3.000 ;
        RECT  8.425 2.740 9.780 3.000 ;
        RECT  8.165 2.295 8.425 3.000 ;
        RECT  6.495 2.740 8.165 3.000 ;
        RECT  6.235 2.620 6.495 3.000 ;
        RECT  5.395 2.740 6.235 3.000 ;
        RECT  5.135 2.620 5.395 3.000 ;
        RECT  2.065 2.740 5.135 3.000 ;
        RECT  1.465 2.570 2.065 3.000 ;
        RECT  0.845 2.740 1.465 3.000 ;
        RECT  0.245 2.365 0.845 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.240 1.230 10.420 1.490 ;
        RECT  10.080 1.230 10.240 2.235 ;
        RECT  9.920 1.230 10.080 1.490 ;
        RECT  9.600 2.075 10.080 2.235 ;
        RECT  9.655 1.735 9.855 1.895 ;
        RECT  9.655 0.765 9.710 1.025 ;
        RECT  9.495 0.765 9.655 1.895 ;
        RECT  9.440 2.075 9.600 2.455 ;
        RECT  9.440 1.135 9.495 1.395 ;
        RECT  8.775 2.295 9.440 2.455 ;
        RECT  9.100 0.745 9.260 2.115 ;
        RECT  8.785 0.745 9.100 0.905 ;
        RECT  8.955 1.855 9.100 2.115 ;
        RECT  8.625 0.310 8.785 0.905 ;
        RECT  8.615 1.955 8.775 2.455 ;
        RECT  7.615 0.310 8.625 0.470 ;
        RECT  8.395 1.955 8.615 2.115 ;
        RECT  8.235 0.650 8.395 2.115 ;
        RECT  7.795 0.650 8.235 0.810 ;
        RECT  7.610 1.955 8.235 2.115 ;
        RECT  7.795 1.470 8.055 1.775 ;
        RECT  7.275 1.470 7.795 1.630 ;
        RECT  7.455 0.310 7.615 1.145 ;
        RECT  7.450 1.815 7.610 2.115 ;
        RECT  6.740 0.310 7.455 0.470 ;
        RECT  7.255 1.815 7.450 1.975 ;
        RECT  7.115 0.650 7.275 1.630 ;
        RECT  6.915 2.185 7.175 2.440 ;
        RECT  7.015 0.650 7.115 0.810 ;
        RECT  7.075 1.470 7.115 1.630 ;
        RECT  6.915 1.470 7.075 1.980 ;
        RECT  6.735 1.720 6.915 1.980 ;
        RECT  4.955 2.280 6.915 2.440 ;
        RECT  6.645 0.990 6.905 1.225 ;
        RECT  6.580 0.310 6.740 0.810 ;
        RECT  6.575 1.720 6.735 2.100 ;
        RECT  6.115 0.990 6.645 1.150 ;
        RECT  4.920 0.650 6.580 0.810 ;
        RECT  5.245 1.940 6.575 2.100 ;
        RECT  5.515 0.990 6.115 1.760 ;
        RECT  4.605 0.990 5.515 1.150 ;
        RECT  5.085 1.455 5.245 2.100 ;
        RECT  4.795 2.280 4.955 2.560 ;
        RECT  4.760 0.365 4.920 0.810 ;
        RECT  4.255 2.400 4.795 2.560 ;
        RECT  3.580 0.650 4.760 0.810 ;
        RECT  4.445 0.990 4.605 2.210 ;
        RECT  3.240 0.310 4.455 0.470 ;
        RECT  4.095 1.165 4.255 2.560 ;
        RECT  3.920 1.165 4.095 1.325 ;
        RECT  2.525 2.400 4.095 2.560 ;
        RECT  3.760 1.065 3.920 1.325 ;
        RECT  3.580 1.545 3.895 1.805 ;
        RECT  3.420 0.650 3.580 2.220 ;
        RECT  2.865 2.060 3.420 2.220 ;
        RECT  3.080 0.310 3.240 1.880 ;
        RECT  3.045 0.430 3.080 0.690 ;
        RECT  3.045 1.620 3.080 1.880 ;
        RECT  2.705 1.600 2.865 2.220 ;
        RECT  1.960 1.600 2.705 1.760 ;
        RECT  2.365 2.055 2.525 2.560 ;
        RECT  1.695 2.055 2.365 2.215 ;
        RECT  1.020 0.310 2.125 0.470 ;
        RECT  1.800 0.680 1.960 1.760 ;
        RECT  1.665 0.680 1.800 0.840 ;
        RECT  1.475 1.600 1.800 1.760 ;
        RECT  1.435 2.055 1.695 2.270 ;
        RECT  1.315 1.470 1.475 1.760 ;
        RECT  1.105 2.055 1.435 2.215 ;
        RECT  1.205 0.650 1.365 1.280 ;
        RECT  1.105 1.120 1.205 1.280 ;
        RECT  0.945 1.120 1.105 2.215 ;
        RECT  0.860 0.310 1.020 0.925 ;
        RECT  0.355 0.765 0.860 0.925 ;
        RECT  0.330 0.765 0.355 1.025 ;
        RECT  0.330 1.790 0.355 2.050 ;
        RECT  0.170 0.765 0.330 2.050 ;
    END
END DFFRHQX8MTH

MACRO DFFRQX1MTH
    CLASS CORE ;
    FOREIGN DFFRQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.915 1.205 8.120 1.365 ;
        RECT  7.755 0.430 7.915 1.365 ;
        RECT  6.695 0.430 7.755 0.590 ;
        RECT  6.535 0.310 6.695 0.590 ;
        RECT  5.340 0.310 6.535 0.470 ;
        RECT  5.180 0.310 5.340 1.150 ;
        RECT  4.475 0.990 5.180 1.150 ;
        RECT  4.315 0.310 4.475 1.150 ;
        RECT  3.070 0.310 4.315 0.470 ;
        RECT  2.910 0.310 3.070 0.640 ;
        RECT  2.390 0.480 2.910 0.640 ;
        RECT  2.230 0.310 2.390 0.640 ;
        RECT  0.750 0.310 2.230 0.470 ;
        RECT  0.590 0.310 0.750 0.760 ;
        RECT  0.360 0.470 0.590 0.760 ;
        RECT  0.200 0.470 0.360 0.870 ;
        END
        AntennaGateArea 0.13 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.730 0.720 8.920 2.145 ;
        RECT  8.705 0.720 8.730 1.170 ;
        RECT  8.635 1.885 8.730 2.145 ;
        RECT  8.635 0.720 8.705 0.980 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.280 1.170 1.785 ;
        END
        AntennaGateArea 0.078 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 0.820 2.810 1.155 ;
        END
        AntennaGateArea 0.0533 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 -0.130 9.020 0.130 ;
        RECT  8.095 -0.130 8.355 0.980 ;
        RECT  7.530 -0.130 8.095 0.130 ;
        RECT  6.930 -0.130 7.530 0.250 ;
        RECT  4.995 -0.130 6.930 0.130 ;
        RECT  4.770 -0.130 4.995 0.810 ;
        RECT  2.730 -0.130 4.770 0.130 ;
        RECT  2.570 -0.130 2.730 0.300 ;
        RECT  0.400 -0.130 2.570 0.130 ;
        RECT  0.140 -0.130 0.400 0.250 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.815 2.740 9.020 3.000 ;
        RECT  8.215 2.570 8.815 3.000 ;
        RECT  7.300 2.740 8.215 3.000 ;
        RECT  7.040 2.570 7.300 3.000 ;
        RECT  5.270 2.740 7.040 3.000 ;
        RECT  5.110 2.245 5.270 3.000 ;
        RECT  0.835 2.740 5.110 3.000 ;
        RECT  0.265 2.360 0.835 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.320 1.265 8.550 1.705 ;
        RECT  8.035 1.545 8.320 1.705 ;
        RECT  7.875 1.545 8.035 2.470 ;
        RECT  7.440 1.545 7.875 1.705 ;
        RECT  7.630 2.225 7.875 2.470 ;
        RECT  6.570 1.885 7.695 2.045 ;
        RECT  7.180 0.865 7.440 1.705 ;
        RECT  6.790 1.325 7.180 1.705 ;
        RECT  5.610 2.385 6.770 2.545 ;
        RECT  6.310 1.885 6.570 2.175 ;
        RECT  6.305 1.885 6.310 2.045 ;
        RECT  6.145 0.650 6.305 2.045 ;
        RECT  6.040 0.650 6.145 0.895 ;
        RECT  5.790 1.330 5.950 2.175 ;
        RECT  5.680 1.330 5.790 1.490 ;
        RECT  5.520 0.685 5.680 1.490 ;
        RECT  5.450 1.670 5.610 2.545 ;
        RECT  4.310 1.330 5.520 1.490 ;
        RECT  4.125 1.670 5.450 1.830 ;
        RECT  3.785 2.010 4.945 2.170 ;
        RECT  3.965 0.650 4.125 1.830 ;
        RECT  3.410 0.650 3.965 0.810 ;
        RECT  3.775 0.990 3.785 2.170 ;
        RECT  3.615 0.990 3.775 2.560 ;
        RECT  1.780 2.400 3.615 2.560 ;
        RECT  3.250 0.650 3.410 2.220 ;
        RECT  2.995 0.820 3.250 1.075 ;
        RECT  3.055 1.675 3.250 2.220 ;
        RECT  1.695 1.675 3.055 1.835 ;
        RECT  2.050 1.335 2.980 1.495 ;
        RECT  2.030 2.015 2.290 2.220 ;
        RECT  1.890 0.695 2.050 1.495 ;
        RECT  1.515 2.015 2.030 2.175 ;
        RECT  1.515 1.010 1.890 1.270 ;
        RECT  1.520 2.355 1.780 2.560 ;
        RECT  1.175 0.650 1.590 0.810 ;
        RECT  1.175 2.400 1.520 2.560 ;
        RECT  1.355 1.010 1.515 2.175 ;
        RECT  1.015 0.650 1.175 1.100 ;
        RECT  1.015 1.965 1.175 2.560 ;
        RECT  0.700 0.940 1.015 1.100 ;
        RECT  0.700 1.965 1.015 2.125 ;
        RECT  0.540 0.940 0.700 2.125 ;
        RECT  0.125 1.895 0.540 2.125 ;
    END
END DFFRQX1MTH

MACRO DFFRQX2MTH
    CLASS CORE ;
    FOREIGN DFFRQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.910 1.205 8.010 1.365 ;
        RECT  7.750 0.430 7.910 1.365 ;
        RECT  6.695 0.430 7.750 0.590 ;
        RECT  6.535 0.310 6.695 0.590 ;
        RECT  5.340 0.310 6.535 0.470 ;
        RECT  5.180 0.310 5.340 1.150 ;
        RECT  4.475 0.990 5.180 1.150 ;
        RECT  4.315 0.310 4.475 1.150 ;
        RECT  3.070 0.310 4.315 0.470 ;
        RECT  2.910 0.310 3.070 0.640 ;
        RECT  2.390 0.480 2.910 0.640 ;
        RECT  2.230 0.310 2.390 0.640 ;
        RECT  0.750 0.310 2.230 0.470 ;
        RECT  0.590 0.310 0.750 0.760 ;
        RECT  0.360 0.470 0.590 0.760 ;
        RECT  0.200 0.470 0.360 0.870 ;
        END
        AntennaGateArea 0.1417 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.380 8.920 2.455 ;
        RECT  8.635 0.380 8.710 0.980 ;
        RECT  8.635 1.855 8.710 2.455 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.280 1.170 1.785 ;
        END
        AntennaGateArea 0.078 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 0.820 2.810 1.155 ;
        END
        AntennaGateArea 0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 -0.130 9.020 0.130 ;
        RECT  8.095 -0.130 8.355 0.980 ;
        RECT  7.530 -0.130 8.095 0.130 ;
        RECT  6.930 -0.130 7.530 0.250 ;
        RECT  4.995 -0.130 6.930 0.130 ;
        RECT  4.770 -0.130 4.995 0.810 ;
        RECT  2.730 -0.130 4.770 0.130 ;
        RECT  2.570 -0.130 2.730 0.300 ;
        RECT  0.400 -0.130 2.570 0.130 ;
        RECT  0.140 -0.130 0.400 0.250 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.295 2.740 9.020 3.000 ;
        RECT  7.035 2.570 7.295 3.000 ;
        RECT  5.290 2.740 7.035 3.000 ;
        RECT  5.130 2.245 5.290 3.000 ;
        RECT  0.835 2.740 5.130 3.000 ;
        RECT  0.265 2.360 0.835 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.370 1.260 8.530 1.705 ;
        RECT  8.030 1.545 8.370 1.705 ;
        RECT  7.870 1.545 8.030 2.470 ;
        RECT  7.320 1.545 7.870 1.705 ;
        RECT  7.630 2.225 7.870 2.470 ;
        RECT  6.530 1.885 7.690 2.045 ;
        RECT  7.060 0.815 7.320 1.705 ;
        RECT  6.790 1.345 7.060 1.705 ;
        RECT  5.630 2.385 6.730 2.545 ;
        RECT  6.310 1.885 6.530 2.175 ;
        RECT  6.270 0.650 6.310 2.175 ;
        RECT  6.150 0.650 6.270 2.045 ;
        RECT  6.040 0.650 6.150 0.895 ;
        RECT  5.810 1.330 5.970 2.175 ;
        RECT  5.680 1.330 5.810 1.490 ;
        RECT  5.520 0.685 5.680 1.490 ;
        RECT  5.470 1.670 5.630 2.545 ;
        RECT  4.310 1.330 5.520 1.490 ;
        RECT  4.125 1.670 5.470 1.830 ;
        RECT  3.780 2.010 4.950 2.170 ;
        RECT  3.965 0.650 4.125 1.830 ;
        RECT  3.410 0.650 3.965 0.810 ;
        RECT  3.620 0.990 3.780 2.560 ;
        RECT  1.780 2.400 3.620 2.560 ;
        RECT  3.250 0.650 3.410 2.220 ;
        RECT  2.995 0.820 3.250 0.980 ;
        RECT  3.060 1.675 3.250 2.220 ;
        RECT  1.695 1.675 3.060 1.835 ;
        RECT  2.050 1.335 2.980 1.495 ;
        RECT  2.030 2.015 2.290 2.220 ;
        RECT  1.890 0.695 2.050 1.495 ;
        RECT  1.515 2.015 2.030 2.175 ;
        RECT  1.625 1.010 1.890 1.170 ;
        RECT  1.520 2.355 1.780 2.560 ;
        RECT  1.515 1.010 1.625 1.270 ;
        RECT  1.175 0.650 1.590 0.810 ;
        RECT  1.175 2.400 1.520 2.560 ;
        RECT  1.355 1.010 1.515 2.175 ;
        RECT  1.015 0.650 1.175 1.100 ;
        RECT  1.015 1.965 1.175 2.560 ;
        RECT  0.700 0.940 1.015 1.100 ;
        RECT  0.700 1.965 1.015 2.125 ;
        RECT  0.540 0.940 0.700 2.125 ;
        RECT  0.125 1.835 0.540 2.125 ;
    END
END DFFRQX2MTH

MACRO DFFRQX4MTH
    CLASS CORE ;
    FOREIGN DFFRQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.845 1.205 8.100 1.365 ;
        RECT  7.685 0.430 7.845 1.365 ;
        RECT  6.695 0.430 7.685 0.590 ;
        RECT  6.535 0.310 6.695 0.590 ;
        RECT  5.340 0.310 6.535 0.470 ;
        RECT  5.180 0.310 5.340 1.150 ;
        RECT  4.475 0.990 5.180 1.150 ;
        RECT  4.315 0.310 4.475 1.150 ;
        RECT  3.070 0.310 4.315 0.470 ;
        RECT  2.910 0.310 3.070 0.640 ;
        RECT  2.390 0.480 2.910 0.640 ;
        RECT  2.230 0.310 2.390 0.640 ;
        RECT  0.750 0.310 2.230 0.470 ;
        RECT  0.590 0.310 0.750 0.760 ;
        RECT  0.360 0.470 0.590 0.760 ;
        RECT  0.200 0.470 0.360 0.870 ;
        END
        AntennaGateArea 0.1794 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.915 1.225 8.985 1.605 ;
        RECT  8.710 0.380 8.915 2.485 ;
        RECT  8.535 0.380 8.710 0.980 ;
        RECT  8.535 1.885 8.710 2.485 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.280 1.170 1.785 ;
        END
        AntennaGateArea 0.078 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 0.820 2.810 1.155 ;
        END
        AntennaGateArea 0.0624 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 -0.130 9.430 0.130 ;
        RECT  9.095 -0.130 9.305 0.985 ;
        RECT  8.285 -0.130 9.095 0.130 ;
        RECT  8.025 -0.130 8.285 0.835 ;
        RECT  7.190 -0.130 8.025 0.130 ;
        RECT  6.930 -0.130 7.190 0.250 ;
        RECT  4.995 -0.130 6.930 0.130 ;
        RECT  4.770 -0.130 4.995 0.810 ;
        RECT  2.730 -0.130 4.770 0.130 ;
        RECT  2.570 -0.130 2.730 0.300 ;
        RECT  0.400 -0.130 2.570 0.130 ;
        RECT  0.140 -0.130 0.400 0.250 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 2.740 9.430 3.000 ;
        RECT  9.095 1.855 9.305 3.000 ;
        RECT  7.295 2.740 9.095 3.000 ;
        RECT  7.035 2.570 7.295 3.000 ;
        RECT  5.290 2.740 7.035 3.000 ;
        RECT  5.130 2.245 5.290 3.000 ;
        RECT  0.835 2.740 5.130 3.000 ;
        RECT  0.265 2.360 0.835 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.370 1.230 8.530 1.705 ;
        RECT  8.030 1.545 8.370 1.705 ;
        RECT  7.870 1.545 8.030 2.470 ;
        RECT  7.450 1.545 7.870 1.705 ;
        RECT  7.585 2.225 7.870 2.470 ;
        RECT  6.530 1.885 7.675 2.045 ;
        RECT  7.190 0.815 7.450 1.705 ;
        RECT  6.790 1.345 7.190 1.705 ;
        RECT  5.630 2.385 6.730 2.545 ;
        RECT  6.310 1.885 6.530 2.175 ;
        RECT  6.270 0.650 6.310 2.175 ;
        RECT  6.150 0.650 6.270 2.045 ;
        RECT  6.040 0.650 6.150 0.895 ;
        RECT  5.810 1.330 5.970 2.175 ;
        RECT  5.680 1.330 5.810 1.490 ;
        RECT  5.520 0.685 5.680 1.490 ;
        RECT  5.470 1.670 5.630 2.545 ;
        RECT  4.310 1.330 5.520 1.490 ;
        RECT  4.125 1.670 5.470 1.830 ;
        RECT  3.780 2.010 4.950 2.170 ;
        RECT  3.965 0.650 4.125 1.830 ;
        RECT  3.410 0.650 3.965 0.810 ;
        RECT  3.620 0.990 3.780 2.560 ;
        RECT  1.780 2.400 3.620 2.560 ;
        RECT  3.250 0.650 3.410 2.220 ;
        RECT  2.995 0.820 3.250 0.980 ;
        RECT  3.060 1.675 3.250 2.220 ;
        RECT  1.695 1.675 3.060 1.835 ;
        RECT  2.050 1.335 2.980 1.495 ;
        RECT  2.030 2.015 2.290 2.220 ;
        RECT  1.890 0.695 2.050 1.495 ;
        RECT  1.515 2.015 2.030 2.175 ;
        RECT  1.625 1.010 1.890 1.170 ;
        RECT  1.520 2.355 1.780 2.560 ;
        RECT  1.515 1.010 1.625 1.270 ;
        RECT  1.175 0.650 1.590 0.810 ;
        RECT  1.175 2.400 1.520 2.560 ;
        RECT  1.355 1.010 1.515 2.175 ;
        RECT  1.015 0.650 1.175 1.100 ;
        RECT  1.015 1.965 1.175 2.560 ;
        RECT  0.700 0.940 1.015 1.100 ;
        RECT  0.700 1.965 1.015 2.125 ;
        RECT  0.540 0.940 0.700 2.125 ;
        RECT  0.125 1.825 0.540 2.125 ;
    END
END DFFRQX4MTH

MACRO DFFRX1MTH
    CLASS CORE ;
    FOREIGN DFFRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.535 1.020 7.120 1.180 ;
        RECT  6.375 0.310 6.535 1.180 ;
        RECT  4.745 0.310 6.375 0.470 ;
        RECT  4.485 0.310 4.745 0.525 ;
        RECT  1.540 0.310 4.485 0.470 ;
        RECT  1.470 0.310 1.540 0.760 ;
        RECT  1.310 0.310 1.470 1.100 ;
        END
        AntennaGateArea 0.13 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 0.815 8.510 1.170 ;
        RECT  8.040 0.815 8.300 1.950 ;
        END
        AntennaDiffArea 0.313 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 0.750 9.330 2.105 ;
        RECT  9.090 0.750 9.170 1.010 ;
        RECT  9.040 1.700 9.170 2.105 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 1.260 0.785 1.640 ;
        END
        AntennaGateArea 0.0767 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.325 2.400 1.735 ;
        RECT  2.010 1.325 2.100 1.545 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.190 -0.130 9.430 0.130 ;
        RECT  8.250 -0.130 9.190 0.295 ;
        RECT  7.690 -0.130 8.250 0.130 ;
        RECT  6.750 -0.130 7.690 0.295 ;
        RECT  0.000 -0.130 6.750 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.585 2.740 9.430 3.000 ;
        RECT  7.985 2.570 8.585 3.000 ;
        RECT  6.905 2.740 7.985 3.000 ;
        RECT  6.645 2.485 6.905 3.000 ;
        RECT  4.295 2.740 6.645 3.000 ;
        RECT  4.035 2.295 4.295 3.000 ;
        RECT  0.000 2.740 4.035 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.910 1.220 8.970 1.480 ;
        RECT  8.750 0.475 8.910 1.480 ;
        RECT  7.750 0.475 8.750 0.635 ;
        RECT  7.675 1.225 7.835 2.305 ;
        RECT  7.590 0.475 7.750 1.010 ;
        RECT  6.860 2.145 7.675 2.305 ;
        RECT  7.465 0.850 7.590 1.010 ;
        RECT  7.305 0.850 7.465 1.965 ;
        RECT  6.805 1.450 7.305 1.610 ;
        RECT  6.700 1.965 6.860 2.305 ;
        RECT  6.545 1.450 6.805 1.710 ;
        RECT  6.195 1.965 6.700 2.125 ;
        RECT  5.745 2.400 6.335 2.560 ;
        RECT  6.035 0.650 6.195 2.125 ;
        RECT  5.855 0.650 6.035 0.810 ;
        RECT  5.925 1.865 6.035 2.125 ;
        RECT  5.745 1.020 5.855 1.180 ;
        RECT  5.585 1.020 5.745 2.560 ;
        RECT  5.060 2.400 5.585 2.560 ;
        RECT  5.405 0.650 5.540 0.810 ;
        RECT  5.245 0.650 5.405 2.125 ;
        RECT  4.165 1.275 5.245 1.435 ;
        RECT  4.900 1.615 5.060 2.560 ;
        RECT  3.895 1.615 4.900 1.775 ;
        RECT  4.475 1.955 4.635 2.395 ;
        RECT  3.525 1.955 4.475 2.115 ;
        RECT  3.735 0.650 3.895 1.775 ;
        RECT  3.165 0.650 3.735 0.810 ;
        RECT  3.365 0.990 3.525 2.115 ;
        RECT  3.355 1.915 3.365 2.115 ;
        RECT  3.195 1.915 3.355 2.560 ;
        RECT  1.075 2.400 3.195 2.560 ;
        RECT  3.005 0.650 3.165 1.735 ;
        RECT  2.825 0.650 3.005 0.810 ;
        RECT  2.845 1.575 3.005 2.220 ;
        RECT  1.455 2.060 2.845 2.220 ;
        RECT  2.620 0.995 2.740 1.395 ;
        RECT  2.580 0.650 2.620 1.395 ;
        RECT  2.460 0.650 2.580 1.155 ;
        RECT  1.940 0.650 2.460 0.810 ;
        RECT  1.810 0.650 1.940 1.150 ;
        RECT  1.810 1.685 1.895 1.845 ;
        RECT  1.780 0.650 1.810 1.845 ;
        RECT  1.650 0.990 1.780 1.845 ;
        RECT  1.635 1.390 1.650 1.845 ;
        RECT  1.130 1.390 1.635 1.550 ;
        RECT  1.295 1.825 1.455 2.220 ;
        RECT  0.695 1.825 1.295 1.985 ;
        RECT  0.970 0.915 1.130 1.550 ;
        RECT  0.915 2.210 1.075 2.560 ;
        RECT  0.600 0.915 0.970 1.075 ;
        RECT  0.260 2.400 0.915 2.560 ;
        RECT  0.440 0.815 0.600 1.075 ;
        RECT  0.260 0.475 0.445 0.635 ;
        RECT  0.100 0.475 0.260 2.560 ;
    END
END DFFRX1MTH

MACRO DFFRX2MTH
    CLASS CORE ;
    FOREIGN DFFRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.320 1.040 7.430 1.200 ;
        RECT  7.160 0.640 7.320 1.200 ;
        RECT  6.700 0.640 7.160 0.800 ;
        RECT  6.540 0.310 6.700 0.800 ;
        RECT  1.540 0.310 6.540 0.470 ;
        RECT  1.325 0.310 1.540 1.100 ;
        END
        AntennaGateArea 0.1417 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.535 0.815 8.635 0.975 ;
        RECT  8.535 1.790 8.635 2.390 ;
        RECT  8.300 0.815 8.535 2.390 ;
        END
        AntennaDiffArea 0.467 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.615 1.700 9.740 2.390 ;
        RECT  9.615 0.400 9.715 1.000 ;
        RECT  9.455 0.400 9.615 2.390 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 1.260 0.805 1.640 ;
        END
        AntennaGateArea 0.0767 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.015 2.360 1.580 ;
        RECT  2.100 1.015 2.150 1.315 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.175 -0.130 9.840 0.130 ;
        RECT  8.915 -0.130 9.175 0.295 ;
        RECT  7.820 -0.130 8.915 0.130 ;
        RECT  7.140 -0.130 7.820 0.300 ;
        RECT  6.880 -0.130 7.140 0.460 ;
        RECT  0.000 -0.130 6.880 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.175 2.740 9.840 3.000 ;
        RECT  8.915 1.790 9.175 3.000 ;
        RECT  7.990 2.740 8.915 3.000 ;
        RECT  7.050 2.465 7.990 3.000 ;
        RECT  4.765 2.740 7.050 3.000 ;
        RECT  4.165 2.285 4.765 3.000 ;
        RECT  0.000 2.740 4.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.115 0.475 9.275 1.480 ;
        RECT  8.060 0.475 9.115 0.635 ;
        RECT  7.900 0.475 8.060 1.540 ;
        RECT  7.575 1.380 7.900 1.540 ;
        RECT  7.235 2.125 7.825 2.285 ;
        RECT  7.415 1.380 7.575 1.945 ;
        RECT  6.880 1.380 7.415 1.540 ;
        RECT  7.075 1.890 7.235 2.285 ;
        RECT  6.270 1.890 7.075 2.050 ;
        RECT  6.720 0.980 6.880 1.540 ;
        RECT  5.820 2.280 6.450 2.440 ;
        RECT  6.110 0.650 6.270 2.050 ;
        RECT  5.985 0.650 6.110 0.810 ;
        RECT  6.005 1.790 6.110 2.050 ;
        RECT  5.820 1.050 5.925 1.210 ;
        RECT  5.660 1.050 5.820 2.440 ;
        RECT  5.105 2.280 5.660 2.440 ;
        RECT  5.480 0.680 5.650 0.840 ;
        RECT  5.320 0.680 5.480 2.050 ;
        RECT  4.190 1.220 5.320 1.380 ;
        RECT  4.945 1.560 5.105 2.440 ;
        RECT  3.920 1.560 4.945 1.720 ;
        RECT  3.550 1.900 4.715 2.060 ;
        RECT  3.760 0.650 3.920 1.720 ;
        RECT  3.040 0.650 3.760 0.810 ;
        RECT  3.400 0.990 3.550 2.060 ;
        RECT  3.390 0.990 3.400 2.555 ;
        RECT  3.240 1.900 3.390 2.555 ;
        RECT  1.075 2.395 3.240 2.555 ;
        RECT  2.880 0.650 3.040 2.210 ;
        RECT  1.415 2.050 2.880 2.210 ;
        RECT  2.540 0.650 2.700 1.800 ;
        RECT  1.910 0.650 2.540 0.810 ;
        RECT  1.910 1.645 1.960 1.805 ;
        RECT  1.750 0.650 1.910 1.805 ;
        RECT  1.700 1.300 1.750 1.805 ;
        RECT  1.145 1.300 1.700 1.460 ;
        RECT  1.255 1.825 1.415 2.210 ;
        RECT  0.665 1.825 1.255 1.985 ;
        RECT  0.985 0.915 1.145 1.460 ;
        RECT  0.915 2.185 1.075 2.555 ;
        RECT  0.600 0.915 0.985 1.075 ;
        RECT  0.260 2.185 0.915 2.345 ;
        RECT  0.440 0.815 0.600 1.075 ;
        RECT  0.260 0.475 0.445 0.635 ;
        RECT  0.100 0.475 0.260 2.345 ;
    END
END DFFRX2MTH

MACRO DFFRX4MTH
    CLASS CORE ;
    FOREIGN DFFRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.320 1.040 7.415 1.200 ;
        RECT  7.155 0.640 7.320 1.200 ;
        RECT  6.730 0.640 7.155 0.800 ;
        RECT  6.570 0.310 6.730 0.800 ;
        RECT  1.540 0.310 6.570 0.470 ;
        RECT  1.330 0.310 1.540 1.100 ;
        END
        AntennaGateArea 0.1794 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.740 0.815 9.005 2.390 ;
        RECT  8.710 0.815 8.740 1.170 ;
        END
        AntennaDiffArea 0.604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.020 1.290 10.150 1.580 ;
        RECT  9.790 0.375 10.020 2.390 ;
        RECT  9.760 0.375 9.790 1.025 ;
        RECT  9.760 1.790 9.790 2.390 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 1.260 0.810 1.640 ;
        END
        AntennaGateArea 0.0767 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.015 2.360 1.580 ;
        RECT  2.100 1.015 2.150 1.315 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 -0.130 10.660 0.130 ;
        RECT  10.275 -0.130 10.535 1.025 ;
        RECT  8.465 -0.130 10.275 0.130 ;
        RECT  8.205 -0.130 8.465 0.295 ;
        RECT  7.175 -0.130 8.205 0.130 ;
        RECT  6.915 -0.130 7.175 0.460 ;
        RECT  0.000 -0.130 6.915 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 2.740 10.660 3.000 ;
        RECT  10.275 1.865 10.535 3.000 ;
        RECT  9.485 2.740 10.275 3.000 ;
        RECT  9.225 1.790 9.485 3.000 ;
        RECT  8.470 2.740 9.225 3.000 ;
        RECT  8.225 1.760 8.470 3.000 ;
        RECT  7.850 2.740 8.225 3.000 ;
        RECT  7.145 2.465 7.850 3.000 ;
        RECT  6.885 2.060 7.145 3.000 ;
        RECT  4.340 2.740 6.885 3.000 ;
        RECT  4.080 2.285 4.340 3.000 ;
        RECT  0.000 2.740 4.080 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.580 1.220 9.610 1.480 ;
        RECT  9.420 0.475 9.580 1.480 ;
        RECT  8.020 0.475 9.420 0.635 ;
        RECT  7.485 2.125 8.045 2.285 ;
        RECT  7.860 0.475 8.020 1.540 ;
        RECT  7.825 1.380 7.860 1.540 ;
        RECT  7.665 1.380 7.825 1.945 ;
        RECT  6.880 1.380 7.665 1.540 ;
        RECT  7.325 1.720 7.485 2.285 ;
        RECT  6.270 1.720 7.325 1.880 ;
        RECT  6.720 0.980 6.880 1.540 ;
        RECT  5.820 2.275 6.450 2.435 ;
        RECT  6.165 0.650 6.270 1.880 ;
        RECT  6.110 0.650 6.165 2.050 ;
        RECT  5.985 0.650 6.110 0.810 ;
        RECT  6.005 1.720 6.110 2.050 ;
        RECT  5.820 1.050 5.920 1.210 ;
        RECT  5.660 1.050 5.820 2.435 ;
        RECT  5.105 2.275 5.660 2.435 ;
        RECT  5.480 0.680 5.650 0.840 ;
        RECT  5.320 0.680 5.480 2.050 ;
        RECT  4.190 1.250 5.320 1.410 ;
        RECT  4.945 1.595 5.105 2.435 ;
        RECT  3.920 1.595 4.945 1.755 ;
        RECT  4.550 1.940 4.710 2.395 ;
        RECT  3.550 1.940 4.550 2.100 ;
        RECT  3.760 0.650 3.920 1.755 ;
        RECT  3.040 0.650 3.760 0.810 ;
        RECT  3.400 0.990 3.550 2.100 ;
        RECT  3.390 0.990 3.400 2.555 ;
        RECT  3.240 1.915 3.390 2.555 ;
        RECT  1.075 2.395 3.240 2.555 ;
        RECT  2.880 0.650 3.040 2.210 ;
        RECT  1.415 2.050 2.880 2.210 ;
        RECT  2.540 0.650 2.700 1.800 ;
        RECT  1.915 0.650 2.540 0.810 ;
        RECT  1.915 1.685 1.945 1.845 ;
        RECT  1.745 0.650 1.915 1.845 ;
        RECT  1.685 1.320 1.745 1.845 ;
        RECT  1.150 1.320 1.685 1.480 ;
        RECT  1.255 1.825 1.415 2.210 ;
        RECT  0.665 1.825 1.255 1.985 ;
        RECT  0.990 0.915 1.150 1.480 ;
        RECT  0.915 2.185 1.075 2.555 ;
        RECT  0.600 0.915 0.990 1.075 ;
        RECT  0.260 2.185 0.915 2.345 ;
        RECT  0.440 0.815 0.600 1.075 ;
        RECT  0.260 0.475 0.445 0.635 ;
        RECT  0.100 0.475 0.260 2.345 ;
    END
END DFFRX4MTH

MACRO DFFSHQX1MTH
    CLASS CORE ;
    FOREIGN DFFSHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.715 1.100 4.080 1.705 ;
        END
        AntennaGateArea 0.1417 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.105 0.760 11.380 2.335 ;
        END
        AntennaDiffArea 0.34 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.875 2.710 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.195 0.965 1.580 ;
        RECT  0.465 1.195 0.510 1.455 ;
        END
        AntennaGateArea 0.1469 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 -0.130 11.480 0.130 ;
        RECT  10.635 -0.130 10.845 0.965 ;
        RECT  8.860 -0.130 10.635 0.130 ;
        RECT  8.600 -0.130 8.860 0.260 ;
        RECT  2.415 -0.130 8.600 0.130 ;
        RECT  2.255 -0.130 2.415 0.300 ;
        RECT  0.580 -0.130 2.255 0.130 ;
        RECT  0.420 -0.130 0.580 0.300 ;
        RECT  0.000 -0.130 0.420 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.795 2.740 11.480 3.000 ;
        RECT  10.635 1.735 10.795 3.000 ;
        RECT  9.890 2.570 10.635 3.000 ;
        RECT  7.300 2.740 9.890 3.000 ;
        RECT  7.040 2.620 7.300 3.000 ;
        RECT  6.140 2.740 7.040 3.000 ;
        RECT  5.880 2.620 6.140 3.000 ;
        RECT  3.650 2.740 5.880 3.000 ;
        RECT  2.710 2.620 3.650 3.000 ;
        RECT  0.735 2.740 2.710 3.000 ;
        RECT  0.235 2.235 0.735 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.455 1.220 10.825 1.480 ;
        RECT  10.295 0.370 10.455 2.335 ;
        RECT  9.710 0.370 10.295 0.530 ;
        RECT  9.620 2.175 10.295 2.335 ;
        RECT  9.905 0.765 10.115 1.995 ;
        RECT  9.625 1.205 9.905 1.470 ;
        RECT  9.450 0.310 9.710 0.530 ;
        RECT  9.445 0.775 9.635 0.935 ;
        RECT  9.460 2.175 9.620 2.455 ;
        RECT  8.400 2.295 9.460 2.455 ;
        RECT  9.165 0.370 9.450 0.530 ;
        RECT  9.285 0.775 9.445 1.775 ;
        RECT  9.200 1.515 9.285 1.775 ;
        RECT  9.040 1.515 9.200 2.115 ;
        RECT  9.005 0.370 9.165 0.635 ;
        RECT  8.520 1.955 9.040 2.115 ;
        RECT  8.300 0.475 9.005 0.635 ;
        RECT  8.700 0.815 8.860 1.775 ;
        RECT  7.960 0.815 8.700 0.975 ;
        RECT  8.360 1.155 8.520 2.115 ;
        RECT  7.620 1.155 8.360 1.315 ;
        RECT  8.140 0.375 8.300 0.635 ;
        RECT  8.020 1.495 8.180 2.440 ;
        RECT  6.680 2.280 8.020 2.440 ;
        RECT  7.800 0.310 7.960 0.975 ;
        RECT  7.720 1.940 7.840 2.100 ;
        RECT  2.755 0.310 7.800 0.470 ;
        RECT  7.560 1.595 7.720 2.100 ;
        RECT  7.460 0.650 7.620 1.315 ;
        RECT  7.280 1.595 7.560 1.755 ;
        RECT  3.535 0.650 7.460 0.810 ;
        RECT  7.120 0.990 7.280 1.755 ;
        RECT  7.020 0.990 7.120 1.150 ;
        RECT  6.360 1.595 7.120 1.755 ;
        RECT  5.550 1.935 6.880 2.095 ;
        RECT  6.580 0.990 6.840 1.415 ;
        RECT  6.420 2.280 6.680 2.500 ;
        RECT  5.550 0.990 6.580 1.150 ;
        RECT  5.570 2.280 6.420 2.440 ;
        RECT  6.100 1.330 6.360 1.755 ;
        RECT  5.410 2.280 5.570 2.490 ;
        RECT  5.390 0.990 5.550 2.095 ;
        RECT  4.890 2.330 5.410 2.490 ;
        RECT  5.230 1.860 5.390 2.095 ;
        RECT  5.070 1.860 5.230 2.120 ;
        RECT  4.890 1.065 4.970 1.325 ;
        RECT  4.730 1.065 4.890 2.490 ;
        RECT  1.585 2.280 4.730 2.440 ;
        RECT  4.390 1.545 4.550 2.100 ;
        RECT  3.050 1.940 4.390 2.100 ;
        RECT  3.375 0.650 3.535 1.760 ;
        RECT  3.230 1.600 3.375 1.760 ;
        RECT  3.095 0.650 3.195 0.810 ;
        RECT  3.050 0.650 3.095 1.420 ;
        RECT  2.935 0.650 3.050 2.100 ;
        RECT  2.890 1.260 2.935 2.100 ;
        RECT  2.720 1.775 2.890 1.935 ;
        RECT  2.595 0.310 2.755 0.665 ;
        RECT  1.850 0.480 2.595 0.665 ;
        RECT  1.850 1.775 2.040 1.935 ;
        RECT  1.685 0.480 1.850 1.935 ;
        RECT  1.515 1.315 1.685 1.575 ;
        RECT  1.335 2.215 1.585 2.500 ;
        RECT  0.920 0.310 1.455 0.470 ;
        RECT  1.175 0.765 1.335 2.500 ;
        RECT  0.760 0.310 0.920 0.930 ;
        RECT  0.385 0.770 0.760 0.930 ;
        RECT  0.285 0.770 0.385 1.025 ;
        RECT  0.285 1.685 0.335 1.945 ;
        RECT  0.125 0.770 0.285 1.945 ;
    END
END DFFSHQX1MTH

MACRO DFFSHQX2MTH
    CLASS CORE ;
    FOREIGN DFFSHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.715 1.100 4.080 1.705 ;
        END
        AntennaGateArea 0.1664 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.105 0.425 11.380 2.335 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.875 2.710 1.485 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.195 0.965 1.580 ;
        RECT  0.465 1.195 0.510 1.455 ;
        END
        AntennaGateArea 0.1599 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 -0.130 11.480 0.130 ;
        RECT  10.635 -0.130 10.845 0.965 ;
        RECT  8.860 -0.130 10.635 0.130 ;
        RECT  8.600 -0.130 8.860 0.260 ;
        RECT  2.415 -0.130 8.600 0.130 ;
        RECT  2.255 -0.130 2.415 0.300 ;
        RECT  0.580 -0.130 2.255 0.130 ;
        RECT  0.420 -0.130 0.580 0.300 ;
        RECT  0.000 -0.130 0.420 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.875 2.740 11.480 3.000 ;
        RECT  10.635 1.735 10.875 3.000 ;
        RECT  9.890 2.570 10.635 3.000 ;
        RECT  7.300 2.740 9.890 3.000 ;
        RECT  7.040 2.620 7.300 3.000 ;
        RECT  6.140 2.740 7.040 3.000 ;
        RECT  5.880 2.620 6.140 3.000 ;
        RECT  3.910 2.740 5.880 3.000 ;
        RECT  3.310 2.620 3.910 3.000 ;
        RECT  2.920 2.740 3.310 3.000 ;
        RECT  2.320 2.620 2.920 3.000 ;
        RECT  0.735 2.740 2.320 3.000 ;
        RECT  0.235 2.235 0.735 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.455 1.220 10.795 1.480 ;
        RECT  10.295 0.380 10.455 2.335 ;
        RECT  9.710 0.380 10.295 0.540 ;
        RECT  9.620 2.175 10.295 2.335 ;
        RECT  9.955 0.765 10.115 1.945 ;
        RECT  9.905 1.205 9.955 1.945 ;
        RECT  9.625 1.205 9.905 1.470 ;
        RECT  9.450 0.355 9.710 0.540 ;
        RECT  9.445 0.775 9.635 0.935 ;
        RECT  9.460 2.175 9.620 2.455 ;
        RECT  8.400 2.295 9.460 2.455 ;
        RECT  9.165 0.380 9.450 0.540 ;
        RECT  9.285 0.775 9.445 1.775 ;
        RECT  9.200 1.515 9.285 1.775 ;
        RECT  9.040 1.515 9.200 2.115 ;
        RECT  9.005 0.380 9.165 0.635 ;
        RECT  8.520 1.955 9.040 2.115 ;
        RECT  8.300 0.475 9.005 0.635 ;
        RECT  8.700 0.815 8.860 1.775 ;
        RECT  7.960 0.815 8.700 0.975 ;
        RECT  8.360 1.155 8.520 2.115 ;
        RECT  7.620 1.155 8.360 1.315 ;
        RECT  8.140 0.375 8.300 0.635 ;
        RECT  8.020 1.495 8.180 2.440 ;
        RECT  6.680 2.280 8.020 2.440 ;
        RECT  7.800 0.310 7.960 0.975 ;
        RECT  7.740 1.940 7.840 2.100 ;
        RECT  2.755 0.310 7.800 0.470 ;
        RECT  7.580 1.595 7.740 2.100 ;
        RECT  7.460 0.650 7.620 1.315 ;
        RECT  7.280 1.595 7.580 1.755 ;
        RECT  3.535 0.650 7.460 0.810 ;
        RECT  7.020 0.990 7.280 1.755 ;
        RECT  6.360 1.595 7.020 1.755 ;
        RECT  5.550 1.935 6.880 2.095 ;
        RECT  6.580 0.990 6.840 1.415 ;
        RECT  6.420 2.280 6.680 2.500 ;
        RECT  5.550 0.990 6.580 1.150 ;
        RECT  5.570 2.280 6.420 2.440 ;
        RECT  6.100 1.330 6.360 1.755 ;
        RECT  5.410 2.280 5.570 2.515 ;
        RECT  5.390 0.990 5.550 2.095 ;
        RECT  4.890 2.355 5.410 2.515 ;
        RECT  5.230 1.915 5.390 2.095 ;
        RECT  5.070 1.915 5.230 2.175 ;
        RECT  4.890 1.065 4.970 1.325 ;
        RECT  4.730 1.065 4.890 2.515 ;
        RECT  1.585 2.280 4.730 2.440 ;
        RECT  4.390 1.545 4.550 2.100 ;
        RECT  3.050 1.940 4.390 2.100 ;
        RECT  3.375 0.650 3.535 1.760 ;
        RECT  3.230 1.600 3.375 1.760 ;
        RECT  3.095 0.650 3.195 0.810 ;
        RECT  3.050 0.650 3.095 1.420 ;
        RECT  2.935 0.650 3.050 2.100 ;
        RECT  2.890 1.260 2.935 2.100 ;
        RECT  2.770 1.685 2.890 2.100 ;
        RECT  2.595 0.310 2.755 0.665 ;
        RECT  1.850 0.480 2.595 0.665 ;
        RECT  1.850 1.735 2.040 1.895 ;
        RECT  1.685 0.480 1.850 1.895 ;
        RECT  1.515 1.315 1.685 1.575 ;
        RECT  1.335 2.235 1.585 2.495 ;
        RECT  0.920 0.310 1.455 0.470 ;
        RECT  1.175 0.765 1.335 2.495 ;
        RECT  0.760 0.310 0.920 0.930 ;
        RECT  0.385 0.770 0.760 0.930 ;
        RECT  0.285 0.770 0.385 1.025 ;
        RECT  0.285 1.685 0.335 1.945 ;
        RECT  0.125 0.770 0.285 1.945 ;
    END
END DFFSHQX2MTH

MACRO DFFSHQX4MTH
    CLASS CORE ;
    FOREIGN DFFSHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.100 4.110 1.705 ;
        END
        AntennaGateArea 0.2002 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.735 1.285 11.790 1.595 ;
        RECT  11.480 0.400 11.735 2.410 ;
        RECT  11.450 0.400 11.480 1.000 ;
        RECT  11.445 1.810 11.480 2.410 ;
        END
        AntennaDiffArea 0.604 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.875 2.705 1.355 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.195 0.885 1.580 ;
        END
        AntennaGateArea 0.2288 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.160 -0.130 12.300 0.130 ;
        RECT  11.920 -0.130 12.160 1.000 ;
        RECT  11.120 -0.130 11.920 0.130 ;
        RECT  10.860 -0.130 11.120 0.250 ;
        RECT  9.300 -0.130 10.860 0.130 ;
        RECT  9.040 -0.130 9.300 0.260 ;
        RECT  2.410 -0.130 9.040 0.130 ;
        RECT  2.250 -0.130 2.410 0.300 ;
        RECT  0.580 -0.130 2.250 0.130 ;
        RECT  0.420 -0.130 0.580 0.300 ;
        RECT  0.000 -0.130 0.420 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.155 2.740 12.300 3.000 ;
        RECT  11.915 1.810 12.155 3.000 ;
        RECT  11.105 2.740 11.915 3.000 ;
        RECT  10.465 2.570 11.105 3.000 ;
        RECT  6.170 2.740 10.465 3.000 ;
        RECT  5.910 2.620 6.170 3.000 ;
        RECT  3.920 2.740 5.910 3.000 ;
        RECT  3.320 2.620 3.920 3.000 ;
        RECT  2.920 2.740 3.320 3.000 ;
        RECT  2.320 2.620 2.920 3.000 ;
        RECT  0.735 2.740 2.320 3.000 ;
        RECT  0.235 2.235 0.735 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.075 1.215 11.275 1.475 ;
        RECT  10.915 0.465 11.075 2.335 ;
        RECT  10.315 0.465 10.915 0.625 ;
        RECT  10.775 1.215 10.915 1.475 ;
        RECT  10.275 2.175 10.915 2.335 ;
        RECT  10.565 1.685 10.665 1.945 ;
        RECT  10.565 0.815 10.615 0.975 ;
        RECT  10.405 0.815 10.565 1.945 ;
        RECT  10.355 0.815 10.405 0.975 ;
        RECT  10.295 1.205 10.405 1.465 ;
        RECT  10.155 0.370 10.315 0.625 ;
        RECT  10.115 2.175 10.275 2.455 ;
        RECT  9.605 0.370 10.155 0.565 ;
        RECT  9.070 2.295 10.115 2.455 ;
        RECT  9.930 1.515 10.025 1.775 ;
        RECT  9.930 0.775 9.985 0.935 ;
        RECT  9.765 0.775 9.930 2.115 ;
        RECT  9.725 0.775 9.765 0.935 ;
        RECT  9.155 1.955 9.765 2.115 ;
        RECT  9.445 0.370 9.605 0.635 ;
        RECT  9.335 0.815 9.495 1.775 ;
        RECT  8.680 0.475 9.445 0.635 ;
        RECT  8.000 0.815 9.335 0.975 ;
        RECT  8.995 1.155 9.155 2.115 ;
        RECT  7.650 1.155 8.995 1.315 ;
        RECT  8.625 1.545 8.785 2.440 ;
        RECT  8.180 0.375 8.680 0.635 ;
        RECT  8.200 1.545 8.625 1.705 ;
        RECT  6.710 2.280 8.625 2.440 ;
        RECT  7.310 1.940 8.445 2.100 ;
        RECT  7.840 0.310 8.000 0.975 ;
        RECT  2.755 0.310 7.840 0.470 ;
        RECT  7.490 0.650 7.650 1.315 ;
        RECT  3.600 0.650 7.490 0.810 ;
        RECT  7.150 0.990 7.310 2.100 ;
        RECT  7.050 0.990 7.150 1.150 ;
        RECT  6.390 1.595 7.150 1.755 ;
        RECT  5.580 1.935 6.910 2.095 ;
        RECT  6.610 0.990 6.870 1.415 ;
        RECT  6.450 2.280 6.710 2.500 ;
        RECT  5.580 0.990 6.610 1.150 ;
        RECT  5.600 2.280 6.450 2.440 ;
        RECT  6.130 1.330 6.390 1.755 ;
        RECT  5.440 2.280 5.600 2.490 ;
        RECT  5.420 0.990 5.580 2.095 ;
        RECT  4.900 2.330 5.440 2.490 ;
        RECT  5.240 1.840 5.420 2.095 ;
        RECT  5.080 1.840 5.240 2.120 ;
        RECT  4.900 1.180 5.000 1.440 ;
        RECT  4.740 1.180 4.900 2.490 ;
        RECT  1.635 2.280 4.740 2.440 ;
        RECT  4.400 1.660 4.560 2.100 ;
        RECT  3.045 1.940 4.400 2.100 ;
        RECT  3.440 0.650 3.600 1.760 ;
        RECT  3.230 1.600 3.440 1.760 ;
        RECT  3.095 0.650 3.195 0.810 ;
        RECT  3.045 0.650 3.095 1.370 ;
        RECT  2.935 0.650 3.045 2.100 ;
        RECT  2.885 1.210 2.935 2.100 ;
        RECT  2.770 1.565 2.885 2.100 ;
        RECT  2.595 0.310 2.755 0.685 ;
        RECT  1.875 0.525 2.595 0.685 ;
        RECT  1.875 1.735 2.040 1.895 ;
        RECT  1.710 0.525 1.875 1.895 ;
        RECT  1.455 1.310 1.710 1.570 ;
        RECT  1.275 2.195 1.635 2.440 ;
        RECT  0.920 0.310 1.525 0.470 ;
        RECT  1.115 0.700 1.275 2.440 ;
        RECT  0.760 0.310 0.920 0.910 ;
        RECT  0.385 0.700 0.760 0.910 ;
        RECT  0.285 0.700 0.385 0.960 ;
        RECT  0.285 1.685 0.335 1.945 ;
        RECT  0.125 0.700 0.285 1.945 ;
    END
END DFFSHQX4MTH

MACRO DFFSHQX8MTH
    CLASS CORE ;
    FOREIGN DFFSHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.100 4.110 1.705 ;
        END
        AntennaGateArea 0.2002 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.635 0.400 12.895 2.370 ;
        RECT  11.890 1.285 12.635 1.595 ;
        RECT  11.595 0.400 11.890 2.410 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.875 2.705 1.355 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.245 0.885 1.580 ;
        END
        AntennaGateArea 0.2288 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 -0.130 13.530 0.130 ;
        RECT  13.145 -0.130 13.405 1.000 ;
        RECT  12.385 -0.130 13.145 0.130 ;
        RECT  12.125 -0.130 12.385 1.000 ;
        RECT  11.415 -0.130 12.125 0.130 ;
        RECT  11.155 -0.130 11.415 1.000 ;
        RECT  10.735 -0.130 11.155 0.270 ;
        RECT  9.315 -0.130 10.735 0.130 ;
        RECT  9.055 -0.130 9.315 0.260 ;
        RECT  2.410 -0.130 9.055 0.130 ;
        RECT  2.180 -0.130 2.410 0.300 ;
        RECT  0.580 -0.130 2.180 0.130 ;
        RECT  0.420 -0.130 0.580 0.300 ;
        RECT  0.000 -0.130 0.420 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.805 13.405 3.000 ;
        RECT  12.385 2.740 13.145 3.000 ;
        RECT  12.125 1.795 12.385 3.000 ;
        RECT  11.325 2.740 12.125 3.000 ;
        RECT  10.385 2.500 11.325 3.000 ;
        RECT  6.170 2.740 10.385 3.000 ;
        RECT  5.910 2.620 6.170 3.000 ;
        RECT  3.920 2.740 5.910 3.000 ;
        RECT  3.320 2.620 3.920 3.000 ;
        RECT  2.920 2.740 3.320 3.000 ;
        RECT  2.320 2.620 2.920 3.000 ;
        RECT  0.735 2.740 2.320 3.000 ;
        RECT  0.235 2.235 0.735 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.055 1.215 11.390 1.475 ;
        RECT  10.975 1.215 11.055 2.285 ;
        RECT  10.895 0.465 10.975 2.285 ;
        RECT  10.815 0.465 10.895 1.475 ;
        RECT  10.205 2.125 10.895 2.285 ;
        RECT  10.315 0.465 10.815 0.625 ;
        RECT  10.635 1.685 10.715 1.945 ;
        RECT  10.375 0.815 10.635 1.945 ;
        RECT  10.295 1.205 10.375 1.465 ;
        RECT  10.155 0.405 10.315 0.625 ;
        RECT  10.045 2.125 10.205 2.455 ;
        RECT  9.585 0.405 10.155 0.565 ;
        RECT  9.070 2.295 10.045 2.455 ;
        RECT  9.865 1.515 10.025 1.775 ;
        RECT  9.865 0.775 9.985 0.935 ;
        RECT  9.700 0.775 9.865 2.115 ;
        RECT  9.155 1.955 9.700 2.115 ;
        RECT  9.425 0.405 9.585 0.635 ;
        RECT  9.335 0.815 9.495 1.775 ;
        RECT  8.680 0.475 9.425 0.635 ;
        RECT  8.000 0.815 9.335 0.975 ;
        RECT  8.995 1.155 9.155 2.115 ;
        RECT  7.650 1.155 8.995 1.315 ;
        RECT  8.610 1.545 8.770 2.440 ;
        RECT  8.180 0.375 8.680 0.635 ;
        RECT  8.200 1.545 8.610 1.705 ;
        RECT  6.710 2.280 8.610 2.440 ;
        RECT  7.310 1.940 8.430 2.100 ;
        RECT  7.840 0.310 8.000 0.975 ;
        RECT  2.755 0.310 7.840 0.470 ;
        RECT  7.490 0.650 7.650 1.315 ;
        RECT  3.600 0.650 7.490 0.810 ;
        RECT  7.150 0.990 7.310 2.100 ;
        RECT  7.050 0.990 7.150 1.150 ;
        RECT  6.390 1.595 7.150 1.755 ;
        RECT  5.660 1.935 6.910 2.095 ;
        RECT  6.610 0.990 6.870 1.415 ;
        RECT  6.450 2.280 6.710 2.500 ;
        RECT  5.660 0.990 6.610 1.150 ;
        RECT  5.600 2.280 6.450 2.440 ;
        RECT  6.130 1.330 6.390 1.755 ;
        RECT  5.500 0.990 5.660 2.095 ;
        RECT  5.440 2.280 5.600 2.500 ;
        RECT  5.420 0.990 5.500 1.150 ;
        RECT  5.240 1.840 5.500 2.095 ;
        RECT  4.900 2.330 5.440 2.500 ;
        RECT  5.080 1.840 5.240 2.120 ;
        RECT  4.900 1.180 5.000 1.440 ;
        RECT  4.740 1.180 4.900 2.500 ;
        RECT  1.635 2.280 4.740 2.440 ;
        RECT  4.400 1.660 4.560 2.100 ;
        RECT  3.045 1.940 4.400 2.100 ;
        RECT  3.440 0.650 3.600 1.760 ;
        RECT  3.230 1.600 3.440 1.760 ;
        RECT  3.095 0.650 3.195 0.810 ;
        RECT  3.045 0.650 3.095 1.370 ;
        RECT  2.935 0.650 3.045 2.100 ;
        RECT  2.885 1.210 2.935 2.100 ;
        RECT  2.770 1.565 2.885 2.100 ;
        RECT  2.595 0.310 2.755 0.685 ;
        RECT  1.875 0.525 2.595 0.685 ;
        RECT  1.875 1.735 2.040 1.895 ;
        RECT  1.710 0.525 1.875 1.895 ;
        RECT  1.455 1.310 1.710 1.570 ;
        RECT  1.275 2.195 1.635 2.440 ;
        RECT  0.920 0.310 1.525 0.470 ;
        RECT  1.115 0.700 1.275 2.440 ;
        RECT  0.760 0.310 0.920 0.910 ;
        RECT  0.285 0.750 0.760 0.910 ;
        RECT  0.285 1.685 0.335 1.945 ;
        RECT  0.125 0.750 0.285 1.945 ;
    END
END DFFSHQX8MTH

MACRO DFFSQX1MTH
    CLASS CORE ;
    FOREIGN DFFSQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.715 1.330 7.420 1.540 ;
        RECT  6.555 1.330 6.715 2.560 ;
        RECT  6.155 2.400 6.555 2.560 ;
        END
        AntennaGateArea 0.1079 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 1.700 8.920 1.990 ;
        RECT  8.735 0.400 8.895 2.390 ;
        RECT  8.635 0.400 8.735 0.660 ;
        RECT  8.710 1.700 8.735 2.390 ;
        RECT  8.635 1.790 8.710 2.390 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 0.880 0.760 1.450 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.320 2.765 1.480 ;
        RECT  1.975 1.320 2.400 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 -0.130 9.020 0.130 ;
        RECT  8.095 -0.130 8.355 0.250 ;
        RECT  7.765 -0.130 8.095 0.130 ;
        RECT  7.165 -0.130 7.765 0.250 ;
        RECT  2.395 -0.130 7.165 0.130 ;
        RECT  2.135 -0.130 2.395 0.250 ;
        RECT  0.725 -0.130 2.135 0.130 ;
        RECT  0.385 -0.130 0.725 0.300 ;
        RECT  0.125 -0.130 0.385 0.640 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.740 9.020 3.000 ;
        RECT  7.755 2.570 8.355 3.000 ;
        RECT  7.475 2.740 7.755 3.000 ;
        RECT  7.215 2.570 7.475 3.000 ;
        RECT  5.975 2.740 7.215 3.000 ;
        RECT  5.375 2.620 5.975 3.000 ;
        RECT  5.185 2.740 5.375 3.000 ;
        RECT  4.585 2.620 5.185 3.000 ;
        RECT  3.740 2.740 4.585 3.000 ;
        RECT  3.580 2.570 3.740 3.000 ;
        RECT  0.410 2.740 3.580 3.000 ;
        RECT  0.150 1.960 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.320 1.190 8.555 1.450 ;
        RECT  8.160 0.605 8.320 2.180 ;
        RECT  7.670 0.605 8.160 0.765 ;
        RECT  7.055 2.020 8.160 2.180 ;
        RECT  7.880 1.265 7.980 1.525 ;
        RECT  7.720 0.990 7.880 1.525 ;
        RECT  5.945 0.990 7.720 1.150 ;
        RECT  6.895 2.020 7.055 2.355 ;
        RECT  6.785 0.605 6.885 0.765 ;
        RECT  6.625 0.310 6.785 0.765 ;
        RECT  3.475 0.310 6.625 0.470 ;
        RECT  5.945 1.880 6.370 2.145 ;
        RECT  5.785 0.765 5.945 2.440 ;
        RECT  4.790 2.280 5.785 2.440 ;
        RECT  5.285 1.910 5.410 2.070 ;
        RECT  5.285 0.650 5.375 1.025 ;
        RECT  5.125 0.650 5.285 2.070 ;
        RECT  4.215 0.650 5.125 0.810 ;
        RECT  4.835 1.310 4.895 1.570 ;
        RECT  4.575 0.990 4.835 1.570 ;
        RECT  4.630 1.990 4.790 2.440 ;
        RECT  4.330 1.410 4.575 1.570 ;
        RECT  4.235 1.410 4.330 2.250 ;
        RECT  4.170 1.410 4.235 2.390 ;
        RECT  4.055 0.650 4.215 1.015 ;
        RECT  4.070 1.990 4.170 2.390 ;
        RECT  3.400 2.230 4.070 2.390 ;
        RECT  3.375 0.800 4.055 0.965 ;
        RECT  3.815 1.190 3.975 1.450 ;
        RECT  3.720 1.290 3.815 1.450 ;
        RECT  3.560 1.290 3.720 1.880 ;
        RECT  2.835 1.720 3.560 1.880 ;
        RECT  3.215 0.310 3.475 0.620 ;
        RECT  3.240 2.230 3.400 2.560 ;
        RECT  3.215 0.800 3.375 1.540 ;
        RECT  0.830 2.400 3.240 2.560 ;
        RECT  2.285 0.800 3.215 0.960 ;
        RECT  3.085 1.380 3.215 1.540 ;
        RECT  1.240 2.060 3.060 2.220 ;
        RECT  2.705 0.410 2.965 0.600 ;
        RECT  2.575 1.690 2.835 1.880 ;
        RECT  1.790 0.440 2.705 0.600 ;
        RECT  1.775 1.720 2.575 1.880 ;
        RECT  2.125 0.800 2.285 1.140 ;
        RECT  2.025 0.980 2.125 1.140 ;
        RECT  1.775 0.310 1.790 0.600 ;
        RECT  1.615 0.310 1.775 1.880 ;
        RECT  1.525 0.310 1.615 0.600 ;
        RECT  1.420 1.520 1.615 1.780 ;
        RECT  1.275 0.770 1.435 1.030 ;
        RECT  1.240 0.870 1.275 1.030 ;
        RECT  1.080 0.870 1.240 2.220 ;
    END
END DFFSQX1MTH

MACRO DFFSQX2MTH
    CLASS CORE ;
    FOREIGN DFFSQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.715 1.330 7.420 1.540 ;
        RECT  6.555 1.330 6.715 2.560 ;
        RECT  6.155 2.400 6.555 2.560 ;
        END
        AntennaGateArea 0.1079 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.735 0.400 8.920 2.390 ;
        RECT  8.635 0.400 8.735 1.000 ;
        RECT  8.635 1.700 8.735 2.390 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.340 1.160 0.760 1.690 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.320 2.765 1.480 ;
        RECT  1.975 1.320 2.400 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 -0.130 9.020 0.130 ;
        RECT  8.095 -0.130 8.355 0.250 ;
        RECT  7.765 -0.130 8.095 0.130 ;
        RECT  7.165 -0.130 7.765 0.250 ;
        RECT  2.395 -0.130 7.165 0.130 ;
        RECT  2.135 -0.130 2.395 0.250 ;
        RECT  0.725 -0.130 2.135 0.130 ;
        RECT  0.385 -0.130 0.725 0.300 ;
        RECT  0.125 -0.130 0.385 0.640 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 2.740 9.020 3.000 ;
        RECT  7.755 2.570 8.355 3.000 ;
        RECT  7.475 2.740 7.755 3.000 ;
        RECT  7.215 2.570 7.475 3.000 ;
        RECT  5.975 2.740 7.215 3.000 ;
        RECT  5.375 2.620 5.975 3.000 ;
        RECT  5.185 2.740 5.375 3.000 ;
        RECT  4.585 2.620 5.185 3.000 ;
        RECT  3.740 2.740 4.585 3.000 ;
        RECT  3.580 2.570 3.740 3.000 ;
        RECT  0.410 2.740 3.580 3.000 ;
        RECT  0.150 1.960 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.320 1.190 8.555 1.450 ;
        RECT  8.160 0.605 8.320 2.180 ;
        RECT  7.670 0.605 8.160 0.765 ;
        RECT  7.055 2.020 8.160 2.180 ;
        RECT  7.880 1.265 7.980 1.525 ;
        RECT  7.720 0.990 7.880 1.525 ;
        RECT  5.945 0.990 7.720 1.150 ;
        RECT  6.895 2.020 7.055 2.355 ;
        RECT  6.785 0.605 6.885 0.765 ;
        RECT  6.625 0.310 6.785 0.765 ;
        RECT  3.475 0.310 6.625 0.470 ;
        RECT  5.945 1.880 6.370 2.145 ;
        RECT  5.785 0.765 5.945 2.440 ;
        RECT  4.790 2.280 5.785 2.440 ;
        RECT  5.285 1.910 5.410 2.070 ;
        RECT  5.285 0.650 5.375 1.025 ;
        RECT  5.125 0.650 5.285 2.070 ;
        RECT  4.215 0.650 5.125 0.810 ;
        RECT  4.835 1.310 4.895 1.570 ;
        RECT  4.575 0.990 4.835 1.570 ;
        RECT  4.630 1.990 4.790 2.440 ;
        RECT  4.330 1.410 4.575 1.570 ;
        RECT  4.235 1.410 4.330 2.250 ;
        RECT  4.170 1.410 4.235 2.390 ;
        RECT  4.055 0.650 4.215 1.015 ;
        RECT  4.070 1.990 4.170 2.390 ;
        RECT  3.400 2.230 4.070 2.390 ;
        RECT  3.375 0.800 4.055 0.965 ;
        RECT  3.815 1.190 3.975 1.450 ;
        RECT  3.720 1.290 3.815 1.450 ;
        RECT  3.560 1.290 3.720 1.880 ;
        RECT  2.835 1.720 3.560 1.880 ;
        RECT  3.215 0.310 3.475 0.620 ;
        RECT  3.240 2.230 3.400 2.560 ;
        RECT  3.215 0.800 3.375 1.540 ;
        RECT  0.830 2.400 3.240 2.560 ;
        RECT  2.285 0.800 3.215 0.960 ;
        RECT  3.085 1.380 3.215 1.540 ;
        RECT  1.240 2.060 3.060 2.220 ;
        RECT  2.705 0.410 2.965 0.600 ;
        RECT  2.575 1.690 2.835 1.880 ;
        RECT  1.790 0.440 2.705 0.600 ;
        RECT  1.775 1.720 2.575 1.880 ;
        RECT  2.125 0.800 2.285 1.140 ;
        RECT  2.025 0.980 2.125 1.140 ;
        RECT  1.775 0.310 1.790 0.600 ;
        RECT  1.615 0.310 1.775 1.880 ;
        RECT  1.525 0.310 1.615 0.600 ;
        RECT  1.420 1.520 1.615 1.780 ;
        RECT  1.275 0.770 1.435 1.030 ;
        RECT  1.240 0.870 1.275 1.030 ;
        RECT  1.080 0.870 1.240 2.220 ;
    END
END DFFSQX2MTH

MACRO DFFSQX4MTH
    CLASS CORE ;
    FOREIGN DFFSQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.690 1.330 7.395 1.540 ;
        RECT  6.530 1.330 6.690 2.560 ;
        RECT  6.130 2.400 6.530 2.560 ;
        END
        AntennaGateArea 0.1079 ;
    END SN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.865 1.700 8.920 1.990 ;
        RECT  8.815 1.700 8.865 2.390 ;
        RECT  8.605 0.400 8.815 2.390 ;
        RECT  8.575 1.790 8.605 2.390 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 1.110 0.735 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.320 2.740 1.480 ;
        RECT  1.950 1.320 2.400 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.275 -0.130 9.430 0.130 ;
        RECT  8.015 -0.130 8.275 0.295 ;
        RECT  7.740 -0.130 8.015 0.130 ;
        RECT  7.140 -0.130 7.740 0.250 ;
        RECT  2.370 -0.130 7.140 0.130 ;
        RECT  2.110 -0.130 2.370 0.250 ;
        RECT  0.725 -0.130 2.110 0.130 ;
        RECT  0.385 -0.130 0.725 0.300 ;
        RECT  0.125 -0.130 0.385 0.640 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 2.740 9.430 3.000 ;
        RECT  9.045 2.170 9.305 3.000 ;
        RECT  8.195 2.740 9.045 3.000 ;
        RECT  7.695 2.570 8.195 3.000 ;
        RECT  7.450 2.740 7.695 3.000 ;
        RECT  7.190 2.570 7.450 3.000 ;
        RECT  5.950 2.740 7.190 3.000 ;
        RECT  5.350 2.620 5.950 3.000 ;
        RECT  5.160 2.740 5.350 3.000 ;
        RECT  4.560 2.620 5.160 3.000 ;
        RECT  3.715 2.740 4.560 3.000 ;
        RECT  3.555 2.570 3.715 3.000 ;
        RECT  0.385 2.740 3.555 3.000 ;
        RECT  0.125 2.140 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.295 1.190 8.425 1.450 ;
        RECT  8.135 0.615 8.295 2.180 ;
        RECT  7.645 0.615 8.135 0.775 ;
        RECT  7.030 2.020 8.135 2.180 ;
        RECT  7.855 1.265 7.955 1.525 ;
        RECT  7.695 0.990 7.855 1.525 ;
        RECT  5.920 0.990 7.695 1.150 ;
        RECT  6.870 2.020 7.030 2.355 ;
        RECT  6.760 0.605 6.860 0.765 ;
        RECT  6.600 0.310 6.760 0.765 ;
        RECT  3.450 0.310 6.600 0.470 ;
        RECT  5.920 1.880 6.345 2.145 ;
        RECT  5.760 0.765 5.920 2.440 ;
        RECT  4.765 2.280 5.760 2.440 ;
        RECT  5.260 1.910 5.385 2.070 ;
        RECT  5.260 0.650 5.350 1.025 ;
        RECT  5.100 0.650 5.260 2.070 ;
        RECT  4.190 0.650 5.100 0.810 ;
        RECT  4.810 1.310 4.870 1.570 ;
        RECT  4.550 0.990 4.810 1.570 ;
        RECT  4.605 1.990 4.765 2.440 ;
        RECT  4.305 1.410 4.550 1.570 ;
        RECT  4.210 1.410 4.305 2.250 ;
        RECT  4.145 1.410 4.210 2.390 ;
        RECT  4.030 0.650 4.190 1.015 ;
        RECT  4.045 1.990 4.145 2.390 ;
        RECT  3.375 2.230 4.045 2.390 ;
        RECT  3.350 0.800 4.030 0.965 ;
        RECT  3.790 1.190 3.950 1.450 ;
        RECT  3.695 1.290 3.790 1.450 ;
        RECT  3.535 1.290 3.695 1.880 ;
        RECT  2.810 1.720 3.535 1.880 ;
        RECT  3.190 0.310 3.450 0.620 ;
        RECT  3.215 2.230 3.375 2.560 ;
        RECT  3.190 0.800 3.350 1.540 ;
        RECT  0.805 2.400 3.215 2.560 ;
        RECT  2.260 0.800 3.190 0.960 ;
        RECT  3.060 1.380 3.190 1.540 ;
        RECT  1.215 2.060 3.035 2.220 ;
        RECT  2.680 0.410 2.940 0.600 ;
        RECT  2.550 1.690 2.810 1.880 ;
        RECT  1.765 0.440 2.680 0.600 ;
        RECT  1.750 1.720 2.550 1.880 ;
        RECT  2.100 0.800 2.260 1.140 ;
        RECT  2.000 0.980 2.100 1.140 ;
        RECT  1.750 0.310 1.765 0.600 ;
        RECT  1.590 0.310 1.750 1.880 ;
        RECT  1.500 0.310 1.590 0.600 ;
        RECT  1.395 1.520 1.590 1.780 ;
        RECT  1.250 0.770 1.410 1.030 ;
        RECT  1.215 0.870 1.250 1.030 ;
        RECT  1.055 0.870 1.215 2.220 ;
    END
END DFFSQX4MTH

MACRO DFFSRHQX1MTH
    CLASS CORE ;
    FOREIGN DFFSRHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.700 1.150 4.000 1.660 ;
        END
        AntennaGateArea 0.1365 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.770 1.385 10.030 1.590 ;
        RECT  7.730 1.430 9.770 1.590 ;
        RECT  7.440 1.330 7.730 1.590 ;
        END
        AntennaGateArea 0.1391 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.220 0.765 13.430 2.115 ;
        RECT  13.145 0.765 13.220 1.025 ;
        RECT  13.145 1.850 13.220 2.115 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.055 2.810 1.540 ;
        END
        AntennaGateArea 0.0598 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.230 0.760 1.860 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.865 -0.130 13.530 0.130 ;
        RECT  12.265 -0.130 12.865 0.295 ;
        RECT  2.410 -0.130 12.265 0.130 ;
        RECT  2.150 -0.130 2.410 0.250 ;
        RECT  0.955 -0.130 2.150 0.130 ;
        RECT  0.695 -0.130 0.955 0.250 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.810 2.740 13.530 3.000 ;
        RECT  12.210 2.570 12.810 3.000 ;
        RECT  7.990 2.740 12.210 3.000 ;
        RECT  7.730 2.620 7.990 3.000 ;
        RECT  7.050 2.740 7.730 3.000 ;
        RECT  6.790 2.620 7.050 3.000 ;
        RECT  5.930 2.740 6.790 3.000 ;
        RECT  5.670 2.620 5.930 3.000 ;
        RECT  4.445 2.740 5.670 3.000 ;
        RECT  4.185 2.620 4.445 3.000 ;
        RECT  2.550 2.740 4.185 3.000 ;
        RECT  2.290 2.620 2.550 3.000 ;
        RECT  0.815 2.740 2.290 3.000 ;
        RECT  0.555 2.620 0.815 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.820 1.200 12.920 1.460 ;
        RECT  12.660 0.475 12.820 2.285 ;
        RECT  11.960 0.475 12.660 0.635 ;
        RECT  11.860 2.125 12.660 2.285 ;
        RECT  12.210 0.815 12.370 1.945 ;
        RECT  11.895 0.815 12.210 0.975 ;
        RECT  11.840 1.195 12.210 1.455 ;
        RECT  11.775 0.355 11.960 0.635 ;
        RECT  11.700 2.125 11.860 2.455 ;
        RECT  9.230 0.355 11.775 0.515 ;
        RECT  11.215 2.295 11.700 2.455 ;
        RECT  11.375 1.565 11.520 1.825 ;
        RECT  11.215 0.715 11.375 2.115 ;
        RECT  11.070 0.715 11.215 0.975 ;
        RECT  10.370 1.955 11.215 2.115 ;
        RECT  10.950 2.295 11.215 2.515 ;
        RECT  10.890 1.515 11.035 1.775 ;
        RECT  9.660 2.295 10.950 2.455 ;
        RECT  10.730 0.695 10.890 1.775 ;
        RECT  9.050 0.695 10.730 0.855 ;
        RECT  10.210 1.035 10.370 2.115 ;
        RECT  8.710 1.035 10.210 1.195 ;
        RECT  9.890 1.865 10.210 2.025 ;
        RECT  9.120 1.815 9.380 2.005 ;
        RECT  8.350 1.845 9.120 2.005 ;
        RECT  8.860 2.185 9.120 2.440 ;
        RECT  8.890 0.310 9.050 0.855 ;
        RECT  2.740 0.310 8.890 0.470 ;
        RECT  6.490 2.280 8.860 2.440 ;
        RECT  8.550 0.650 8.710 1.195 ;
        RECT  3.520 0.650 8.550 0.810 ;
        RECT  8.210 0.990 8.370 1.250 ;
        RECT  8.190 1.845 8.350 2.100 ;
        RECT  7.175 0.990 8.210 1.150 ;
        RECT  7.175 1.940 8.190 2.100 ;
        RECT  7.015 0.990 7.175 2.100 ;
        RECT  6.790 0.990 7.015 1.150 ;
        RECT  6.730 1.470 7.015 1.730 ;
        RECT  5.390 0.990 6.590 1.250 ;
        RECT  6.230 2.280 6.490 2.560 ;
        RECT  6.030 1.840 6.290 2.100 ;
        RECT  5.360 2.280 6.230 2.440 ;
        RECT  5.390 1.840 6.030 2.000 ;
        RECT  5.230 0.990 5.390 2.000 ;
        RECT  5.200 2.280 5.360 2.460 ;
        RECT  5.020 1.840 5.230 2.000 ;
        RECT  4.680 2.300 5.200 2.460 ;
        RECT  4.860 1.840 5.020 2.120 ;
        RECT  4.680 1.005 4.930 1.265 ;
        RECT  4.530 1.005 4.680 2.460 ;
        RECT  4.520 1.005 4.530 2.440 ;
        RECT  4.015 2.280 4.520 2.440 ;
        RECT  4.180 1.325 4.340 2.100 ;
        RECT  3.770 1.940 4.180 2.100 ;
        RECT  3.855 2.280 4.015 2.460 ;
        RECT  2.855 2.300 3.855 2.460 ;
        RECT  3.610 1.940 3.770 2.120 ;
        RECT  3.180 1.960 3.610 2.120 ;
        RECT  3.360 0.650 3.520 1.780 ;
        RECT  3.020 0.650 3.180 2.120 ;
        RECT  2.920 0.650 3.020 0.810 ;
        RECT  2.800 1.735 3.020 1.895 ;
        RECT  2.695 2.245 2.855 2.460 ;
        RECT  2.580 0.310 2.740 0.665 ;
        RECT  1.100 2.245 2.695 2.405 ;
        RECT  2.035 0.505 2.580 0.665 ;
        RECT  1.845 0.505 2.035 1.945 ;
        RECT  1.285 1.660 1.845 1.945 ;
        RECT  0.385 0.430 1.655 0.590 ;
        RECT  1.100 0.815 1.525 0.975 ;
        RECT  0.940 0.815 1.100 2.405 ;
        RECT  0.285 0.430 0.385 1.040 ;
        RECT  0.285 2.075 0.385 2.335 ;
        RECT  0.125 0.430 0.285 2.335 ;
    END
END DFFSRHQX1MTH

MACRO DFFSRHQX2MTH
    CLASS CORE ;
    FOREIGN DFFSRHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.700 1.150 4.000 1.660 ;
        END
        AntennaGateArea 0.1586 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.890 1.385 10.150 1.590 ;
        RECT  7.730 1.430 9.890 1.590 ;
        RECT  7.440 1.330 7.730 1.590 ;
        END
        AntennaGateArea 0.1677 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.220 0.380 13.430 2.430 ;
        RECT  13.145 0.380 13.220 0.980 ;
        RECT  13.145 1.830 13.220 2.430 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.055 2.810 1.540 ;
        END
        AntennaGateArea 0.0598 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.210 0.760 1.830 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.865 -0.130 13.530 0.130 ;
        RECT  12.265 -0.130 12.865 0.295 ;
        RECT  2.410 -0.130 12.265 0.130 ;
        RECT  2.150 -0.130 2.410 0.250 ;
        RECT  0.955 -0.130 2.150 0.130 ;
        RECT  0.695 -0.130 0.955 0.250 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.810 2.740 13.530 3.000 ;
        RECT  12.210 2.570 12.810 3.000 ;
        RECT  7.990 2.740 12.210 3.000 ;
        RECT  7.730 2.620 7.990 3.000 ;
        RECT  7.050 2.740 7.730 3.000 ;
        RECT  6.790 2.620 7.050 3.000 ;
        RECT  5.930 2.740 6.790 3.000 ;
        RECT  5.670 2.620 5.930 3.000 ;
        RECT  4.445 2.740 5.670 3.000 ;
        RECT  4.185 2.620 4.445 3.000 ;
        RECT  2.625 2.740 4.185 3.000 ;
        RECT  2.365 2.620 2.625 3.000 ;
        RECT  0.815 2.740 2.365 3.000 ;
        RECT  0.555 2.620 0.815 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.710 1.215 13.035 1.475 ;
        RECT  12.550 0.475 12.710 2.285 ;
        RECT  11.960 0.475 12.550 0.635 ;
        RECT  12.435 1.215 12.550 1.475 ;
        RECT  11.970 2.125 12.550 2.285 ;
        RECT  12.225 1.685 12.370 1.945 ;
        RECT  12.065 0.815 12.225 1.945 ;
        RECT  11.900 0.815 12.065 0.975 ;
        RECT  11.840 1.255 12.065 1.515 ;
        RECT  11.810 2.125 11.970 2.455 ;
        RECT  11.775 0.355 11.960 0.635 ;
        RECT  11.215 2.295 11.810 2.455 ;
        RECT  9.230 0.355 11.775 0.515 ;
        RECT  11.355 0.715 11.515 2.115 ;
        RECT  11.215 0.715 11.355 0.975 ;
        RECT  10.690 1.955 11.355 2.115 ;
        RECT  10.950 2.295 11.215 2.515 ;
        RECT  10.875 0.695 11.035 1.775 ;
        RECT  9.660 2.295 10.950 2.455 ;
        RECT  9.050 0.695 10.875 0.855 ;
        RECT  10.530 1.035 10.690 2.115 ;
        RECT  8.710 1.035 10.530 1.195 ;
        RECT  9.890 1.865 10.530 2.025 ;
        RECT  8.350 1.815 9.380 1.975 ;
        RECT  8.860 2.185 9.120 2.440 ;
        RECT  8.890 0.310 9.050 0.855 ;
        RECT  2.740 0.310 8.890 0.470 ;
        RECT  6.490 2.280 8.860 2.440 ;
        RECT  8.550 0.650 8.710 1.195 ;
        RECT  3.520 0.650 8.550 0.810 ;
        RECT  8.210 0.990 8.370 1.250 ;
        RECT  8.190 1.815 8.350 2.100 ;
        RECT  7.260 0.990 8.210 1.150 ;
        RECT  7.260 1.940 8.190 2.100 ;
        RECT  7.100 0.990 7.260 2.100 ;
        RECT  6.790 0.990 7.100 1.150 ;
        RECT  6.730 1.470 7.100 1.730 ;
        RECT  5.560 0.990 6.590 1.250 ;
        RECT  6.230 2.280 6.490 2.560 ;
        RECT  5.560 1.940 6.290 2.100 ;
        RECT  5.360 2.280 6.230 2.440 ;
        RECT  5.400 0.990 5.560 2.100 ;
        RECT  5.350 0.990 5.400 1.250 ;
        RECT  5.020 1.840 5.400 2.100 ;
        RECT  5.200 2.280 5.360 2.460 ;
        RECT  4.680 2.300 5.200 2.460 ;
        RECT  4.860 1.840 5.020 2.120 ;
        RECT  4.680 1.005 4.930 1.265 ;
        RECT  4.530 1.005 4.680 2.460 ;
        RECT  4.520 1.005 4.530 2.440 ;
        RECT  4.015 2.280 4.520 2.440 ;
        RECT  4.180 1.325 4.340 2.100 ;
        RECT  3.770 1.940 4.180 2.100 ;
        RECT  3.855 2.280 4.015 2.460 ;
        RECT  2.890 2.300 3.855 2.460 ;
        RECT  3.610 1.940 3.770 2.120 ;
        RECT  3.180 1.960 3.610 2.120 ;
        RECT  3.360 0.650 3.520 1.780 ;
        RECT  3.020 0.650 3.180 2.120 ;
        RECT  2.920 0.650 3.020 0.810 ;
        RECT  2.800 1.735 3.020 1.895 ;
        RECT  2.730 2.245 2.890 2.460 ;
        RECT  2.580 0.310 2.740 0.665 ;
        RECT  1.320 2.245 2.730 2.405 ;
        RECT  2.030 0.505 2.580 0.665 ;
        RECT  1.845 0.505 2.030 1.945 ;
        RECT  1.500 1.685 1.845 1.945 ;
        RECT  0.910 0.430 1.655 0.590 ;
        RECT  1.320 0.815 1.525 0.975 ;
        RECT  1.160 0.815 1.320 2.405 ;
        RECT  0.750 0.430 0.910 0.975 ;
        RECT  0.285 0.815 0.750 0.975 ;
        RECT  0.285 2.075 0.385 2.335 ;
        RECT  0.125 0.815 0.285 2.335 ;
    END
END DFFSRHQX2MTH

MACRO DFFSRHQX4MTH
    CLASS CORE ;
    FOREIGN DFFSRHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.155 4.150 1.725 ;
        END
        AntennaGateArea 0.1807 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.185 1.385 10.445 1.635 ;
        RECT  8.970 1.475 10.185 1.635 ;
        RECT  8.710 1.440 8.970 1.635 ;
        RECT  8.140 1.475 8.710 1.635 ;
        RECT  7.850 1.330 8.140 1.635 ;
        RECT  7.670 1.440 7.850 1.635 ;
        END
        AntennaGateArea 0.2041 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.680 1.290 13.840 1.580 ;
        RECT  13.420 0.400 13.680 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.880 2.830 1.580 ;
        END
        AntennaGateArea 0.1313 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.285 1.045 1.675 ;
        END
        AntennaGateArea 0.1807 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 -0.130 14.350 0.130 ;
        RECT  13.965 -0.130 14.225 1.025 ;
        RECT  13.120 -0.130 13.965 0.130 ;
        RECT  12.900 -0.130 13.120 1.005 ;
        RECT  1.650 -0.130 12.900 0.130 ;
        RECT  0.710 -0.130 1.650 0.250 ;
        RECT  0.000 -0.130 0.710 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 2.740 14.350 3.000 ;
        RECT  13.965 1.775 14.225 3.000 ;
        RECT  13.110 2.740 13.965 3.000 ;
        RECT  12.510 2.570 13.110 3.000 ;
        RECT  7.250 2.740 12.510 3.000 ;
        RECT  6.990 2.620 7.250 3.000 ;
        RECT  6.140 2.740 6.990 3.000 ;
        RECT  5.880 2.620 6.140 3.000 ;
        RECT  4.060 2.740 5.880 3.000 ;
        RECT  3.800 2.620 4.060 3.000 ;
        RECT  2.700 2.740 3.800 3.000 ;
        RECT  2.440 2.620 2.700 3.000 ;
        RECT  0.910 2.740 2.440 3.000 ;
        RECT  0.310 2.520 0.910 3.000 ;
        RECT  0.000 2.740 0.310 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.000 1.185 13.165 1.445 ;
        RECT  12.840 1.185 13.000 2.285 ;
        RECT  12.720 1.185 12.840 1.445 ;
        RECT  12.140 2.125 12.840 2.285 ;
        RECT  12.560 0.355 12.720 1.445 ;
        RECT  12.500 1.685 12.660 1.945 ;
        RECT  9.560 0.355 12.560 0.515 ;
        RECT  12.380 1.685 12.500 1.845 ;
        RECT  12.220 0.765 12.380 1.845 ;
        RECT  12.130 1.195 12.220 1.455 ;
        RECT  11.980 2.125 12.140 2.455 ;
        RECT  11.505 2.295 11.980 2.455 ;
        RECT  11.680 1.625 11.860 1.885 ;
        RECT  11.520 0.715 11.680 2.115 ;
        RECT  10.785 1.955 11.520 2.115 ;
        RECT  11.240 2.295 11.505 2.515 ;
        RECT  11.200 1.515 11.330 1.775 ;
        RECT  9.950 2.295 11.240 2.455 ;
        RECT  11.040 0.695 11.200 1.775 ;
        RECT  9.380 0.695 11.040 0.855 ;
        RECT  10.625 1.035 10.785 2.115 ;
        RECT  9.040 1.035 10.625 1.195 ;
        RECT  10.180 1.865 10.625 2.025 ;
        RECT  9.410 1.815 9.670 2.005 ;
        RECT  8.910 1.845 9.410 2.005 ;
        RECT  9.150 2.185 9.410 2.440 ;
        RECT  9.220 0.310 9.380 0.855 ;
        RECT  2.230 0.310 9.220 0.470 ;
        RECT  6.700 2.280 9.150 2.440 ;
        RECT  8.880 0.650 9.040 1.195 ;
        RECT  8.750 1.845 8.910 2.100 ;
        RECT  3.610 0.650 8.880 0.810 ;
        RECT  7.180 1.940 8.750 2.100 ;
        RECT  8.540 0.990 8.700 1.250 ;
        RECT  7.180 0.990 8.540 1.150 ;
        RECT  7.020 0.990 7.180 2.100 ;
        RECT  6.930 1.455 7.020 1.715 ;
        RECT  6.510 1.025 6.840 1.185 ;
        RECT  6.440 2.280 6.700 2.560 ;
        RECT  6.350 1.025 6.510 2.100 ;
        RECT  5.570 2.280 6.440 2.440 ;
        RECT  6.240 1.840 6.350 2.100 ;
        RECT  5.700 1.840 6.240 2.000 ;
        RECT  5.700 0.990 5.750 1.150 ;
        RECT  5.540 0.990 5.700 2.000 ;
        RECT  5.410 2.280 5.570 2.470 ;
        RECT  5.490 0.990 5.540 1.150 ;
        RECT  5.230 1.840 5.540 2.000 ;
        RECT  4.890 2.300 5.410 2.470 ;
        RECT  5.070 1.840 5.230 2.120 ;
        RECT  4.890 1.180 5.020 1.440 ;
        RECT  4.730 1.180 4.890 2.470 ;
        RECT  1.385 2.280 4.730 2.440 ;
        RECT  4.390 1.660 4.550 2.100 ;
        RECT  3.170 1.940 4.390 2.100 ;
        RECT  3.450 0.650 3.610 1.730 ;
        RECT  3.350 1.570 3.450 1.730 ;
        RECT  3.170 0.650 3.270 0.810 ;
        RECT  3.010 0.650 3.170 2.100 ;
        RECT  2.840 1.760 3.010 2.020 ;
        RECT  2.070 0.310 2.230 1.930 ;
        RECT  1.950 0.545 2.070 0.805 ;
        RECT  1.900 1.515 2.070 1.930 ;
        RECT  1.565 1.515 1.900 1.775 ;
        RECT  1.770 1.010 1.885 1.270 ;
        RECT  1.610 0.475 1.770 1.270 ;
        RECT  0.880 0.475 1.610 0.635 ;
        RECT  1.385 0.815 1.415 0.975 ;
        RECT  1.225 0.815 1.385 2.440 ;
        RECT  1.155 0.815 1.225 0.975 ;
        RECT  0.720 0.475 0.880 0.925 ;
        RECT  0.385 0.765 0.720 0.925 ;
        RECT  0.285 0.765 0.385 1.025 ;
        RECT  0.285 1.940 0.385 2.200 ;
        RECT  0.125 0.765 0.285 2.200 ;
    END
END DFFSRHQX4MTH

MACRO DFFSRHQX8MTH
    CLASS CORE ;
    FOREIGN DFFSRHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.090 4.140 1.715 ;
        END
        AntennaGateArea 0.1807 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.185 1.385 10.445 1.635 ;
        RECT  8.140 1.475 10.185 1.635 ;
        RECT  7.915 1.330 8.140 1.635 ;
        RECT  7.850 1.330 7.915 1.600 ;
        RECT  7.670 1.440 7.850 1.600 ;
        END
        AntennaGateArea 0.2041 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.605 0.400 14.865 2.285 ;
        RECT  13.780 1.290 14.605 1.580 ;
        RECT  13.520 0.400 13.780 2.285 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.880 2.830 1.505 ;
        END
        AntennaGateArea 0.1313 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.140 0.760 1.750 ;
        END
        AntennaGateArea 0.1807 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.410 -0.130 15.580 0.130 ;
        RECT  15.150 -0.130 15.410 1.025 ;
        RECT  14.325 -0.130 15.150 0.130 ;
        RECT  14.065 -0.130 14.325 1.025 ;
        RECT  13.120 -0.130 14.065 0.130 ;
        RECT  12.900 -0.130 13.120 1.005 ;
        RECT  0.625 -0.130 12.900 0.130 ;
        RECT  0.365 -0.130 0.625 0.250 ;
        RECT  0.000 -0.130 0.365 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.410 2.740 15.580 3.000 ;
        RECT  15.150 1.755 15.410 3.000 ;
        RECT  14.325 2.740 15.150 3.000 ;
        RECT  14.065 1.760 14.325 3.000 ;
        RECT  13.110 2.740 14.065 3.000 ;
        RECT  12.510 2.570 13.110 3.000 ;
        RECT  7.250 2.740 12.510 3.000 ;
        RECT  6.990 2.620 7.250 3.000 ;
        RECT  6.100 2.740 6.990 3.000 ;
        RECT  5.840 2.620 6.100 3.000 ;
        RECT  4.250 2.740 5.840 3.000 ;
        RECT  3.990 2.620 4.250 3.000 ;
        RECT  2.700 2.740 3.990 3.000 ;
        RECT  2.440 2.620 2.700 3.000 ;
        RECT  0.910 2.740 2.440 3.000 ;
        RECT  0.310 2.520 0.910 3.000 ;
        RECT  0.000 2.740 0.310 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.000 1.185 13.180 1.445 ;
        RECT  12.840 1.185 13.000 2.285 ;
        RECT  12.720 1.185 12.840 1.445 ;
        RECT  12.030 2.125 12.840 2.285 ;
        RECT  12.560 0.475 12.720 1.445 ;
        RECT  12.500 1.685 12.660 1.945 ;
        RECT  12.210 0.475 12.560 0.635 ;
        RECT  12.280 1.685 12.500 1.845 ;
        RECT  12.280 0.815 12.380 0.975 ;
        RECT  12.120 0.815 12.280 1.845 ;
        RECT  12.025 0.355 12.210 0.635 ;
        RECT  11.870 2.125 12.030 2.455 ;
        RECT  9.560 0.355 12.025 0.515 ;
        RECT  11.505 2.295 11.870 2.455 ;
        RECT  11.690 1.565 11.800 1.825 ;
        RECT  11.530 0.715 11.690 2.115 ;
        RECT  10.785 1.955 11.530 2.115 ;
        RECT  11.240 2.295 11.505 2.515 ;
        RECT  11.180 1.515 11.320 1.775 ;
        RECT  9.950 2.295 11.240 2.455 ;
        RECT  11.020 0.695 11.180 1.775 ;
        RECT  9.380 0.695 11.020 0.855 ;
        RECT  10.625 1.035 10.785 2.115 ;
        RECT  9.040 1.035 10.625 1.195 ;
        RECT  10.180 1.865 10.625 2.025 ;
        RECT  9.410 1.815 9.670 2.005 ;
        RECT  8.910 1.845 9.410 2.005 ;
        RECT  9.150 2.185 9.410 2.440 ;
        RECT  9.220 0.310 9.380 0.855 ;
        RECT  2.160 0.310 9.220 0.470 ;
        RECT  6.700 2.280 9.150 2.440 ;
        RECT  8.880 0.650 9.040 1.195 ;
        RECT  8.750 1.845 8.910 2.100 ;
        RECT  3.610 0.650 8.880 0.810 ;
        RECT  7.180 1.940 8.750 2.100 ;
        RECT  8.540 0.990 8.700 1.250 ;
        RECT  7.180 0.990 8.540 1.150 ;
        RECT  7.020 0.990 7.180 2.100 ;
        RECT  6.930 1.455 7.020 1.715 ;
        RECT  6.510 1.025 6.840 1.185 ;
        RECT  6.440 2.280 6.700 2.560 ;
        RECT  6.350 1.025 6.510 2.100 ;
        RECT  5.570 2.280 6.440 2.440 ;
        RECT  6.240 1.840 6.350 2.100 ;
        RECT  5.480 1.840 6.240 2.000 ;
        RECT  5.480 0.990 5.750 1.150 ;
        RECT  5.410 2.280 5.570 2.485 ;
        RECT  5.320 0.990 5.480 2.000 ;
        RECT  4.830 2.300 5.410 2.485 ;
        RECT  5.230 1.840 5.320 2.000 ;
        RECT  5.030 1.840 5.230 2.120 ;
        RECT  4.830 1.180 5.020 1.440 ;
        RECT  4.730 1.180 4.830 2.485 ;
        RECT  4.670 1.180 4.730 2.440 ;
        RECT  1.285 2.280 4.670 2.440 ;
        RECT  4.320 1.485 4.480 2.100 ;
        RECT  3.170 1.940 4.320 2.100 ;
        RECT  3.450 0.650 3.610 1.730 ;
        RECT  3.350 1.570 3.450 1.730 ;
        RECT  3.170 0.650 3.270 0.810 ;
        RECT  3.010 0.650 3.170 2.100 ;
        RECT  2.840 1.695 3.010 1.955 ;
        RECT  2.000 0.310 2.160 1.930 ;
        RECT  1.950 0.550 2.000 0.810 ;
        RECT  1.505 1.570 2.000 1.930 ;
        RECT  1.770 1.035 1.820 1.295 ;
        RECT  1.610 0.310 1.770 1.295 ;
        RECT  0.955 0.310 1.610 0.470 ;
        RECT  1.285 0.650 1.430 0.810 ;
        RECT  1.125 0.650 1.285 2.440 ;
        RECT  0.795 0.310 0.955 0.590 ;
        RECT  0.385 0.430 0.795 0.590 ;
        RECT  0.285 0.430 0.385 0.810 ;
        RECT  0.285 1.945 0.385 2.205 ;
        RECT  0.220 0.430 0.285 2.205 ;
        RECT  0.125 0.650 0.220 2.205 ;
    END
END DFFSRHQX8MTH

MACRO DFFSRX1MTH
    CLASS CORE ;
    FOREIGN DFFSRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.630 1.825 10.890 2.425 ;
        RECT  10.350 2.110 10.630 2.425 ;
        END
        AntennaGateArea 0.1118 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.180 1.330 4.860 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.855 0.735 13.015 1.965 ;
        RECT  12.400 0.735 12.855 0.895 ;
        RECT  12.200 1.805 12.855 1.965 ;
        RECT  12.240 0.635 12.400 0.895 ;
        RECT  11.990 1.805 12.200 2.400 ;
        END
        AntennaDiffArea 0.305 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.195 0.755 13.430 2.125 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.445 1.690 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.110 4.000 1.580 ;
        RECT  3.605 1.110 3.790 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.340 -0.130 13.530 0.130 ;
        RECT  12.740 -0.130 13.340 0.345 ;
        RECT  11.510 -0.130 12.740 0.130 ;
        RECT  11.250 -0.130 11.510 0.345 ;
        RECT  4.380 -0.130 11.250 0.130 ;
        RECT  3.780 -0.130 4.380 0.250 ;
        RECT  2.225 -0.130 3.780 0.130 ;
        RECT  2.065 -0.130 2.225 0.980 ;
        RECT  0.505 -0.130 2.065 0.130 ;
        RECT  0.245 -0.130 0.505 0.965 ;
        RECT  0.000 -0.130 0.245 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.865 2.740 13.530 3.000 ;
        RECT  12.605 2.245 12.865 3.000 ;
        RECT  11.800 2.740 12.605 3.000 ;
        RECT  11.640 1.905 11.800 3.000 ;
        RECT  2.270 2.740 11.640 3.000 ;
        RECT  2.270 2.295 2.320 2.455 ;
        RECT  2.110 2.295 2.270 3.000 ;
        RECT  2.060 2.295 2.110 2.455 ;
        RECT  0.445 2.740 2.110 3.000 ;
        RECT  0.285 2.155 0.445 3.000 ;
        RECT  0.000 2.740 0.285 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.510 1.315 12.670 1.625 ;
        RECT  12.060 1.465 12.510 1.625 ;
        RECT  11.900 0.605 12.060 1.625 ;
        RECT  11.680 0.605 11.900 0.765 ;
        RECT  11.230 1.465 11.900 1.625 ;
        RECT  8.630 1.095 11.650 1.255 ;
        RECT  11.070 1.465 11.230 1.945 ;
        RECT  9.580 1.465 11.070 1.625 ;
        RECT  10.760 0.310 10.920 0.760 ;
        RECT  9.075 0.310 10.760 0.470 ;
        RECT  8.290 0.755 10.280 0.915 ;
        RECT  9.950 2.015 10.050 2.175 ;
        RECT  9.790 2.015 9.950 2.560 ;
        RECT  6.310 2.400 9.790 2.560 ;
        RECT  8.970 1.595 9.310 1.855 ;
        RECT  8.475 0.310 9.075 0.575 ;
        RECT  8.810 1.595 8.970 2.220 ;
        RECT  7.160 2.060 8.810 2.220 ;
        RECT  8.470 1.095 8.630 1.880 ;
        RECT  7.465 0.310 8.475 0.470 ;
        RECT  8.120 1.720 8.470 1.880 ;
        RECT  8.130 0.755 8.290 1.540 ;
        RECT  7.600 1.380 8.130 1.540 ;
        RECT  7.790 0.655 7.950 1.200 ;
        RECT  6.540 1.040 7.790 1.200 ;
        RECT  7.480 1.380 7.600 1.615 ;
        RECT  7.320 1.380 7.480 1.760 ;
        RECT  7.275 0.310 7.465 0.845 ;
        RECT  5.895 1.600 7.320 1.760 ;
        RECT  7.200 0.685 7.275 0.845 ;
        RECT  7.000 1.955 7.160 2.220 ;
        RECT  5.870 1.955 7.000 2.115 ;
        RECT  6.420 1.040 6.540 1.420 ;
        RECT  6.260 0.310 6.420 1.420 ;
        RECT  6.050 2.295 6.310 2.560 ;
        RECT  4.720 0.310 6.260 0.470 ;
        RECT  5.735 0.650 5.895 1.760 ;
        RECT  5.710 1.955 5.870 2.220 ;
        RECT  2.745 2.400 5.840 2.560 ;
        RECT  5.060 0.650 5.735 0.810 ;
        RECT  3.085 2.060 5.710 2.220 ;
        RECT  5.340 0.990 5.530 1.880 ;
        RECT  5.250 0.990 5.340 1.150 ;
        RECT  4.360 1.720 5.340 1.880 ;
        RECT  4.900 0.650 5.060 0.930 ;
        RECT  3.425 0.770 4.900 0.930 ;
        RECT  4.560 0.310 4.720 0.590 ;
        RECT  2.565 0.430 4.560 0.590 ;
        RECT  3.425 1.720 3.645 1.880 ;
        RECT  3.265 0.770 3.425 1.880 ;
        RECT  3.085 1.175 3.265 1.435 ;
        RECT  2.925 1.615 3.085 2.220 ;
        RECT  2.905 0.770 3.035 0.930 ;
        RECT  2.905 1.615 2.925 1.775 ;
        RECT  2.745 0.770 2.905 1.775 ;
        RECT  0.965 1.615 2.745 1.775 ;
        RECT  2.585 1.955 2.745 2.560 ;
        RECT  1.735 1.955 2.585 2.115 ;
        RECT  2.405 0.430 2.565 1.345 ;
        RECT  1.810 1.185 2.405 1.345 ;
        RECT  1.575 1.955 1.735 2.175 ;
        RECT  0.785 2.015 1.575 2.175 ;
        RECT  1.175 0.720 1.335 1.365 ;
        RECT  0.785 1.205 1.175 1.365 ;
        RECT  0.625 1.205 0.785 2.175 ;
    END
END DFFSRX1MTH

MACRO DFFSRX2MTH
    CLASS CORE ;
    FOREIGN DFFSRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.630 1.800 10.890 2.400 ;
        RECT  10.350 2.110 10.630 2.400 ;
        END
        AntennaGateArea 0.1352 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.180 1.330 4.860 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.335 1.685 12.650 1.950 ;
        RECT  12.175 0.765 12.335 1.950 ;
        END
        AntennaDiffArea 0.494 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.195 0.390 13.430 2.400 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.445 1.690 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.110 4.000 1.580 ;
        RECT  3.605 1.110 3.790 1.540 ;
        END
        AntennaGateArea 0.1183 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.895 -0.130 13.530 0.130 ;
        RECT  12.635 -0.130 12.895 0.985 ;
        RECT  4.380 -0.130 12.635 0.130 ;
        RECT  3.780 -0.130 4.380 0.250 ;
        RECT  2.225 -0.130 3.780 0.130 ;
        RECT  2.065 -0.130 2.225 0.995 ;
        RECT  0.505 -0.130 2.065 0.130 ;
        RECT  0.245 -0.130 0.505 0.965 ;
        RECT  0.000 -0.130 0.245 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.865 2.740 13.530 3.000 ;
        RECT  12.605 2.470 12.865 3.000 ;
        RECT  11.845 2.740 12.605 3.000 ;
        RECT  11.585 2.470 11.845 3.000 ;
        RECT  2.270 2.740 11.585 3.000 ;
        RECT  2.270 2.295 2.320 2.455 ;
        RECT  2.110 2.295 2.270 3.000 ;
        RECT  2.060 2.295 2.110 2.455 ;
        RECT  0.445 2.740 2.110 3.000 ;
        RECT  0.285 2.155 0.445 3.000 ;
        RECT  0.000 2.740 0.285 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.855 1.205 13.015 2.290 ;
        RECT  11.995 2.130 12.855 2.290 ;
        RECT  11.835 0.355 11.995 2.290 ;
        RECT  11.680 0.355 11.835 0.515 ;
        RECT  11.230 2.130 11.835 2.290 ;
        RECT  11.495 1.095 11.655 1.420 ;
        RECT  8.630 1.095 11.495 1.255 ;
        RECT  11.070 1.445 11.230 2.290 ;
        RECT  10.200 1.445 11.070 1.605 ;
        RECT  10.710 0.310 10.970 0.760 ;
        RECT  9.075 0.310 10.710 0.470 ;
        RECT  8.290 0.755 10.280 0.915 ;
        RECT  9.580 1.445 10.200 1.635 ;
        RECT  9.950 1.965 10.050 2.225 ;
        RECT  9.790 1.965 9.950 2.560 ;
        RECT  6.310 2.400 9.790 2.560 ;
        RECT  8.970 1.595 9.310 1.855 ;
        RECT  8.475 0.310 9.075 0.575 ;
        RECT  8.810 1.595 8.970 2.220 ;
        RECT  7.160 2.060 8.810 2.220 ;
        RECT  8.470 1.095 8.630 1.880 ;
        RECT  7.460 0.310 8.475 0.470 ;
        RECT  8.120 1.720 8.470 1.880 ;
        RECT  8.130 0.755 8.290 1.540 ;
        RECT  7.600 1.380 8.130 1.540 ;
        RECT  7.790 0.655 7.950 1.200 ;
        RECT  6.540 1.040 7.790 1.200 ;
        RECT  7.480 1.380 7.600 1.615 ;
        RECT  7.320 1.380 7.480 1.760 ;
        RECT  7.200 0.310 7.460 0.835 ;
        RECT  5.895 1.600 7.320 1.760 ;
        RECT  7.000 1.955 7.160 2.220 ;
        RECT  5.870 1.955 7.000 2.115 ;
        RECT  6.420 1.040 6.540 1.420 ;
        RECT  6.260 0.310 6.420 1.420 ;
        RECT  6.050 2.295 6.310 2.560 ;
        RECT  4.720 0.310 6.260 0.470 ;
        RECT  5.735 0.650 5.895 1.760 ;
        RECT  5.710 1.955 5.870 2.220 ;
        RECT  2.745 2.400 5.840 2.560 ;
        RECT  5.060 0.650 5.735 0.810 ;
        RECT  3.085 2.060 5.710 2.220 ;
        RECT  5.340 0.990 5.530 1.880 ;
        RECT  5.250 0.990 5.340 1.150 ;
        RECT  4.360 1.720 5.340 1.880 ;
        RECT  4.900 0.650 5.060 0.930 ;
        RECT  3.425 0.770 4.900 0.930 ;
        RECT  4.560 0.310 4.720 0.590 ;
        RECT  2.565 0.430 4.560 0.590 ;
        RECT  3.425 1.720 3.645 1.880 ;
        RECT  3.265 0.770 3.425 1.880 ;
        RECT  3.085 1.175 3.265 1.435 ;
        RECT  2.925 1.615 3.085 2.220 ;
        RECT  2.905 0.785 3.035 0.945 ;
        RECT  2.905 1.615 2.925 1.775 ;
        RECT  2.745 0.785 2.905 1.775 ;
        RECT  0.965 1.615 2.745 1.775 ;
        RECT  2.585 1.955 2.745 2.560 ;
        RECT  1.735 1.955 2.585 2.115 ;
        RECT  2.405 0.430 2.565 1.345 ;
        RECT  1.805 1.185 2.405 1.345 ;
        RECT  1.575 1.955 1.735 2.175 ;
        RECT  0.785 2.015 1.575 2.175 ;
        RECT  1.175 0.735 1.335 1.365 ;
        RECT  0.785 1.205 1.175 1.365 ;
        RECT  0.625 1.205 0.785 2.175 ;
    END
END DFFSRX2MTH

MACRO DFFSRX4MTH
    CLASS CORE ;
    FOREIGN DFFSRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.325 1.820 10.585 2.420 ;
        RECT  9.940 2.110 10.325 2.420 ;
        END
        AntennaGateArea 0.1521 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 1.330 4.450 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.610 0.390 12.645 0.990 ;
        RECT  12.400 0.390 12.610 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.740 1.290 13.925 1.580 ;
        RECT  13.505 0.425 13.740 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.320 0.355 1.580 ;
        RECT  0.100 0.880 0.310 1.580 ;
        END
        AntennaGateArea 0.0715 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 1.110 3.590 1.580 ;
        RECT  3.305 1.190 3.350 1.450 ;
        END
        AntennaGateArea 0.1443 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 -0.130 14.350 0.130 ;
        RECT  13.965 -0.130 14.225 0.955 ;
        RECT  13.205 -0.130 13.965 0.130 ;
        RECT  12.945 -0.130 13.205 0.955 ;
        RECT  12.155 -0.130 12.945 0.130 ;
        RECT  11.555 -0.130 12.155 0.300 ;
        RECT  11.100 -0.130 11.555 0.130 ;
        RECT  10.810 -0.130 11.100 0.825 ;
        RECT  3.970 -0.130 10.810 0.130 ;
        RECT  3.370 -0.130 3.970 0.250 ;
        RECT  2.930 -0.130 3.370 0.130 ;
        RECT  1.990 -0.130 2.930 0.250 ;
        RECT  0.385 -0.130 1.990 0.130 ;
        RECT  0.125 -0.130 0.385 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 2.740 14.350 3.000 ;
        RECT  13.965 1.865 14.225 3.000 ;
        RECT  13.175 2.740 13.965 3.000 ;
        RECT  12.915 2.525 13.175 3.000 ;
        RECT  12.095 2.740 12.915 3.000 ;
        RECT  11.155 2.570 12.095 3.000 ;
        RECT  1.995 2.740 11.155 3.000 ;
        RECT  1.835 2.245 1.995 3.000 ;
        RECT  1.065 2.740 1.835 3.000 ;
        RECT  0.125 2.620 1.065 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.165 1.285 13.325 2.330 ;
        RECT  12.140 2.170 13.165 2.330 ;
        RECT  11.980 0.750 12.140 2.330 ;
        RECT  11.325 0.750 11.980 0.910 ;
        RECT  11.295 1.735 11.980 1.895 ;
        RECT  11.510 1.095 11.770 1.435 ;
        RECT  8.220 1.095 11.510 1.255 ;
        RECT  11.135 1.465 11.295 1.895 ;
        RECT  9.170 1.465 11.135 1.625 ;
        RECT  10.300 0.310 10.560 0.915 ;
        RECT  8.665 0.310 10.300 0.470 ;
        RECT  7.880 0.755 9.870 0.915 ;
        RECT  9.540 2.015 9.640 2.175 ;
        RECT  9.380 2.015 9.540 2.560 ;
        RECT  5.870 2.400 9.380 2.560 ;
        RECT  8.560 1.595 8.900 1.855 ;
        RECT  8.065 0.310 8.665 0.575 ;
        RECT  8.400 1.595 8.560 2.220 ;
        RECT  6.750 2.060 8.400 2.220 ;
        RECT  8.060 1.095 8.220 1.880 ;
        RECT  7.050 0.310 8.065 0.470 ;
        RECT  7.710 1.720 8.060 1.880 ;
        RECT  7.720 0.755 7.880 1.540 ;
        RECT  7.220 1.380 7.720 1.540 ;
        RECT  7.380 0.655 7.540 1.200 ;
        RECT  6.130 1.040 7.380 1.200 ;
        RECT  7.100 1.380 7.220 1.615 ;
        RECT  6.940 1.380 7.100 1.760 ;
        RECT  6.880 0.310 7.050 0.840 ;
        RECT  5.495 1.600 6.940 1.760 ;
        RECT  6.790 0.680 6.880 0.840 ;
        RECT  6.590 1.955 6.750 2.220 ;
        RECT  5.430 1.955 6.590 2.115 ;
        RECT  6.010 1.040 6.130 1.420 ;
        RECT  5.850 0.310 6.010 1.420 ;
        RECT  5.610 2.295 5.870 2.560 ;
        RECT  4.310 0.310 5.850 0.470 ;
        RECT  5.335 0.650 5.495 1.760 ;
        RECT  5.270 1.955 5.430 2.220 ;
        RECT  2.335 2.400 5.430 2.560 ;
        RECT  4.650 0.650 5.335 0.810 ;
        RECT  2.675 2.060 5.270 2.220 ;
        RECT  4.940 0.990 5.100 1.880 ;
        RECT  4.840 0.990 4.940 1.150 ;
        RECT  3.950 1.720 4.940 1.880 ;
        RECT  4.490 0.650 4.650 0.930 ;
        RECT  3.125 0.770 4.490 0.930 ;
        RECT  4.150 0.310 4.310 0.590 ;
        RECT  1.785 0.430 4.150 0.590 ;
        RECT  3.125 1.720 3.235 1.880 ;
        RECT  2.965 0.770 3.125 1.880 ;
        RECT  2.535 1.110 2.965 1.270 ;
        RECT  2.195 0.770 2.785 0.930 ;
        RECT  2.515 1.565 2.675 2.220 ;
        RECT  2.375 1.110 2.535 1.370 ;
        RECT  2.195 1.565 2.515 1.725 ;
        RECT  2.175 1.905 2.335 2.560 ;
        RECT  2.035 0.770 2.195 1.725 ;
        RECT  1.310 1.905 2.175 2.065 ;
        RECT  1.425 0.770 2.035 0.930 ;
        RECT  1.625 0.330 1.785 0.590 ;
        RECT  1.265 0.310 1.425 0.930 ;
        RECT  1.150 1.230 1.310 2.175 ;
        RECT  0.740 0.310 1.265 0.470 ;
        RECT  1.085 1.230 1.150 1.390 ;
        RECT  0.845 2.015 1.150 2.175 ;
        RECT  0.925 0.725 1.085 1.390 ;
        RECT  0.740 1.575 0.885 1.835 ;
        RECT  0.580 0.310 0.740 1.835 ;
    END
END DFFSRX4MTH

MACRO DFFSX1MTH
    CLASS CORE ;
    FOREIGN DFFSX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.750 1.330 7.320 1.620 ;
        RECT  6.620 1.460 6.750 1.620 ;
        RECT  6.460 1.460 6.620 2.560 ;
        RECT  5.865 2.400 6.460 2.560 ;
        END
        AntennaGateArea 0.1118 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.280 0.865 8.440 1.990 ;
        RECT  8.070 0.865 8.280 1.025 ;
        RECT  7.890 1.700 8.280 1.990 ;
        END
        AntennaDiffArea 0.344 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 0.740 9.330 2.070 ;
        RECT  9.045 0.740 9.170 1.000 ;
        RECT  9.120 1.700 9.170 2.070 ;
        RECT  9.045 1.810 9.120 2.070 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.560 1.700 0.720 1.990 ;
        RECT  0.400 1.355 0.560 1.990 ;
        END
        AntennaGateArea 0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.320 2.755 1.510 ;
        RECT  2.110 1.320 2.400 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.150 -0.130 9.430 0.130 ;
        RECT  8.210 -0.130 9.150 0.250 ;
        RECT  7.390 -0.130 8.210 0.130 ;
        RECT  6.790 -0.130 7.390 0.300 ;
        RECT  2.385 -0.130 6.790 0.130 ;
        RECT  1.785 -0.130 2.385 0.250 ;
        RECT  0.725 -0.130 1.785 0.130 ;
        RECT  0.385 -0.130 0.725 0.300 ;
        RECT  0.125 -0.130 0.385 0.640 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.245 2.740 9.430 3.000 ;
        RECT  6.985 2.620 7.245 3.000 ;
        RECT  5.670 2.740 6.985 3.000 ;
        RECT  4.730 2.620 5.670 3.000 ;
        RECT  0.395 2.740 4.730 3.000 ;
        RECT  0.135 2.175 0.395 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.780 1.190 8.990 1.450 ;
        RECT  8.620 0.435 8.780 2.330 ;
        RECT  7.960 0.435 8.620 0.595 ;
        RECT  6.960 2.170 8.620 2.330 ;
        RECT  7.660 1.315 8.100 1.475 ;
        RECT  7.700 0.355 7.960 0.595 ;
        RECT  7.500 0.990 7.660 1.475 ;
        RECT  6.280 0.990 7.500 1.150 ;
        RECT  6.460 0.640 6.990 0.800 ;
        RECT  6.800 2.170 6.960 2.440 ;
        RECT  6.300 0.310 6.460 0.800 ;
        RECT  3.975 0.310 6.300 0.470 ;
        RECT  6.120 0.990 6.280 2.130 ;
        RECT  5.890 0.815 6.120 1.150 ;
        RECT  6.020 1.930 6.120 2.130 ;
        RECT  5.600 1.970 6.020 2.130 ;
        RECT  5.550 0.865 5.710 1.790 ;
        RECT  5.440 1.970 5.600 2.440 ;
        RECT  5.130 0.865 5.550 1.025 ;
        RECT  5.260 1.630 5.550 1.790 ;
        RECT  4.640 2.280 5.440 2.440 ;
        RECT  4.790 1.210 5.370 1.450 ;
        RECT  5.100 1.630 5.260 2.090 ;
        RECT  4.970 0.650 5.130 1.025 ;
        RECT  5.000 1.930 5.100 2.090 ;
        RECT  4.350 0.650 4.970 0.810 ;
        RECT  4.530 0.990 4.790 1.450 ;
        RECT  4.480 1.880 4.640 2.440 ;
        RECT  4.240 1.290 4.530 1.450 ;
        RECT  4.190 0.650 4.350 0.945 ;
        RECT  4.080 1.290 4.240 2.560 ;
        RECT  3.465 0.785 4.190 0.945 ;
        RECT  3.920 2.135 4.080 2.560 ;
        RECT  3.715 0.310 3.975 0.570 ;
        RECT  0.830 2.400 3.920 2.560 ;
        RECT  3.740 1.510 3.900 1.880 ;
        RECT  2.760 1.720 3.740 1.880 ;
        RECT  3.270 0.410 3.465 0.945 ;
        RECT  3.205 0.410 3.270 1.540 ;
        RECT  3.010 0.785 3.205 1.540 ;
        RECT  2.275 0.785 3.010 0.945 ;
        RECT  1.240 2.060 2.980 2.220 ;
        RECT  2.695 0.360 2.955 0.590 ;
        RECT  2.500 1.690 2.760 1.880 ;
        RECT  1.835 0.430 2.695 0.590 ;
        RECT  1.835 1.720 2.500 1.880 ;
        RECT  2.115 0.785 2.275 1.135 ;
        RECT  2.015 0.975 2.115 1.135 ;
        RECT  1.675 0.430 1.835 1.880 ;
        RECT  1.345 0.430 1.675 0.590 ;
        RECT  1.420 1.590 1.675 1.850 ;
        RECT  1.335 0.770 1.495 1.030 ;
        RECT  1.085 0.335 1.345 0.590 ;
        RECT  1.240 0.870 1.335 1.030 ;
        RECT  1.080 0.870 1.240 2.220 ;
    END
END DFFSX1MTH

MACRO DFFSX2MTH
    CLASS CORE ;
    FOREIGN DFFSX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.750 1.330 7.320 1.620 ;
        RECT  6.590 1.460 6.750 1.620 ;
        RECT  6.430 1.460 6.590 2.560 ;
        RECT  5.830 2.400 6.430 2.560 ;
        END
        AntennaGateArea 0.1352 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.460 0.815 8.630 0.975 ;
        RECT  8.460 1.695 8.570 1.990 ;
        RECT  8.300 0.815 8.460 1.990 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 1.700 9.740 1.990 ;
        RECT  9.425 0.400 9.685 2.390 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.545 1.610 ;
        END
        AntennaGateArea 0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.320 2.755 1.510 ;
        RECT  2.110 1.320 2.400 1.540 ;
        END
        AntennaGateArea 0.1183 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 -0.130 9.840 0.130 ;
        RECT  8.910 -0.130 9.170 0.250 ;
        RECT  8.030 -0.130 8.910 0.130 ;
        RECT  7.430 -0.130 8.030 0.250 ;
        RECT  2.385 -0.130 7.430 0.130 ;
        RECT  1.445 -0.130 2.385 0.250 ;
        RECT  0.795 -0.130 1.445 0.130 ;
        RECT  0.455 -0.130 0.795 0.300 ;
        RECT  0.195 -0.130 0.455 0.640 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.140 2.740 9.840 3.000 ;
        RECT  8.880 2.570 9.140 3.000 ;
        RECT  7.830 2.740 8.880 3.000 ;
        RECT  6.890 2.570 7.830 3.000 ;
        RECT  5.645 2.740 6.890 3.000 ;
        RECT  4.705 2.620 5.645 3.000 ;
        RECT  0.410 2.740 4.705 3.000 ;
        RECT  0.150 1.790 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.060 1.190 9.240 1.450 ;
        RECT  9.030 0.435 9.060 1.450 ;
        RECT  8.870 0.435 9.030 2.375 ;
        RECT  8.120 0.435 8.870 0.595 ;
        RECT  8.090 2.215 8.870 2.375 ;
        RECT  7.860 0.435 8.120 0.810 ;
        RECT  7.830 1.870 8.090 2.375 ;
        RECT  6.930 2.215 7.830 2.375 ;
        RECT  7.625 0.990 7.785 1.525 ;
        RECT  6.250 0.990 7.625 1.150 ;
        RECT  7.050 0.600 7.135 0.760 ;
        RECT  6.875 0.310 7.050 0.760 ;
        RECT  6.770 2.095 6.930 2.375 ;
        RECT  4.035 0.310 6.875 0.470 ;
        RECT  6.090 0.815 6.250 2.130 ;
        RECT  6.030 0.815 6.090 1.075 ;
        RECT  5.990 1.940 6.090 2.130 ;
        RECT  5.580 1.970 5.990 2.130 ;
        RECT  5.585 0.865 5.745 1.790 ;
        RECT  5.430 0.865 5.585 1.025 ;
        RECT  5.230 1.630 5.585 1.790 ;
        RECT  5.420 1.970 5.580 2.440 ;
        RECT  5.270 0.650 5.430 1.025 ;
        RECT  4.640 2.280 5.420 2.440 ;
        RECT  5.035 1.210 5.405 1.450 ;
        RECT  4.465 0.650 5.270 0.810 ;
        RECT  5.070 1.630 5.230 2.100 ;
        RECT  4.970 1.940 5.070 2.100 ;
        RECT  4.775 0.990 5.035 1.450 ;
        RECT  4.240 1.290 4.775 1.450 ;
        RECT  4.480 1.900 4.640 2.440 ;
        RECT  4.305 0.650 4.465 1.110 ;
        RECT  3.465 0.950 4.305 1.110 ;
        RECT  4.080 1.290 4.240 2.560 ;
        RECT  3.920 2.135 4.080 2.560 ;
        RECT  3.775 0.310 4.035 0.520 ;
        RECT  0.830 2.400 3.920 2.560 ;
        RECT  3.740 1.530 3.900 1.880 ;
        RECT  2.760 1.720 3.740 1.880 ;
        RECT  3.270 0.360 3.465 1.110 ;
        RECT  3.205 0.360 3.270 1.540 ;
        RECT  3.010 0.950 3.205 1.540 ;
        RECT  2.150 0.950 3.010 1.110 ;
        RECT  1.240 2.060 2.980 2.220 ;
        RECT  2.695 0.340 2.955 0.590 ;
        RECT  2.500 1.690 2.760 1.880 ;
        RECT  1.710 0.430 2.695 0.590 ;
        RECT  1.710 1.720 2.500 1.880 ;
        RECT  1.890 0.950 2.150 1.140 ;
        RECT  1.550 0.430 1.710 1.880 ;
        RECT  1.235 0.430 1.550 0.590 ;
        RECT  1.420 1.590 1.550 1.880 ;
        RECT  1.240 0.770 1.365 1.030 ;
        RECT  1.205 0.770 1.240 2.220 ;
        RECT  0.975 0.310 1.235 0.590 ;
        RECT  1.080 0.870 1.205 2.220 ;
    END
END DFFSX2MTH

MACRO DFFSX4MTH
    CLASS CORE ;
    FOREIGN DFFSX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.030 1.330 7.320 1.800 ;
        RECT  6.010 1.330 7.030 1.490 ;
        RECT  5.850 1.330 6.010 1.765 ;
        RECT  5.780 1.605 5.850 1.765 ;
        RECT  5.620 1.605 5.780 1.880 ;
        END
        AntennaGateArea 0.2002 ;
    END SN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.785 0.805 8.920 0.965 ;
        RECT  8.605 0.805 8.785 1.955 ;
        RECT  8.260 1.700 8.605 1.955 ;
        END
        AntennaDiffArea 0.608 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.025 1.290 10.150 1.580 ;
        RECT  9.765 0.405 10.025 2.400 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.190 0.460 1.580 ;
        END
        AntennaGateArea 0.0988 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 0.830 2.465 1.130 ;
        END
        AntennaGateArea 0.1482 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.540 -0.130 10.660 0.130 ;
        RECT  10.280 -0.130 10.540 0.990 ;
        RECT  9.465 -0.130 10.280 0.130 ;
        RECT  9.205 -0.130 9.465 0.285 ;
        RECT  8.150 -0.130 9.205 0.130 ;
        RECT  7.550 -0.130 8.150 0.300 ;
        RECT  7.365 -0.130 7.550 0.130 ;
        RECT  7.135 -0.130 7.365 0.810 ;
        RECT  1.890 -0.130 7.135 0.130 ;
        RECT  1.290 -0.130 1.890 0.250 ;
        RECT  0.390 -0.130 1.290 0.130 ;
        RECT  0.130 -0.130 0.390 0.300 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 2.740 10.660 3.000 ;
        RECT  10.275 1.825 10.535 3.000 ;
        RECT  9.505 2.740 10.275 3.000 ;
        RECT  9.305 1.805 9.505 3.000 ;
        RECT  9.170 2.570 9.305 3.000 ;
        RECT  8.290 2.740 9.170 3.000 ;
        RECT  8.030 2.480 8.290 3.000 ;
        RECT  7.080 2.740 8.030 3.000 ;
        RECT  6.820 2.580 7.080 3.000 ;
        RECT  6.220 2.740 6.820 3.000 ;
        RECT  5.620 2.570 6.220 3.000 ;
        RECT  3.520 2.740 5.620 3.000 ;
        RECT  3.320 2.570 3.520 3.000 ;
        RECT  0.390 2.740 3.320 3.000 ;
        RECT  0.130 2.570 0.390 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.260 1.190 9.530 1.450 ;
        RECT  9.125 0.465 9.260 1.450 ;
        RECT  9.100 0.465 9.125 2.295 ;
        RECT  8.425 0.465 9.100 0.625 ;
        RECT  8.965 1.190 9.100 2.295 ;
        RECT  7.730 2.135 8.965 2.295 ;
        RECT  8.265 0.465 8.425 0.775 ;
        RECT  7.710 0.615 8.265 0.775 ;
        RECT  7.715 1.170 8.055 1.430 ;
        RECT  7.470 2.135 7.730 2.430 ;
        RECT  7.555 0.990 7.715 1.430 ;
        RECT  5.810 0.990 7.555 1.150 ;
        RECT  6.795 2.135 7.470 2.295 ;
        RECT  6.720 0.525 6.820 0.785 ;
        RECT  6.635 1.845 6.795 2.295 ;
        RECT  6.560 0.310 6.720 0.785 ;
        RECT  6.535 1.845 6.635 2.005 ;
        RECT  3.450 0.310 6.560 0.470 ;
        RECT  5.855 2.065 6.115 2.265 ;
        RECT  5.440 2.105 5.855 2.265 ;
        RECT  5.670 0.750 5.810 1.150 ;
        RECT  5.510 0.750 5.670 1.395 ;
        RECT  5.440 1.235 5.510 1.395 ;
        RECT  5.280 1.235 5.440 2.560 ;
        RECT  4.585 2.400 5.280 2.560 ;
        RECT  5.100 0.740 5.250 1.000 ;
        RECT  4.940 0.650 5.100 2.220 ;
        RECT  3.940 0.650 4.940 0.810 ;
        RECT  4.835 2.060 4.940 2.220 ;
        RECT  4.670 0.990 4.730 1.150 ;
        RECT  4.520 0.990 4.670 1.520 ;
        RECT  4.325 2.260 4.585 2.560 ;
        RECT  4.360 0.990 4.520 2.080 ;
        RECT  4.025 1.920 4.360 2.080 ;
        RECT  3.650 1.580 4.075 1.740 ;
        RECT  3.865 1.920 4.025 2.390 ;
        RECT  3.730 0.650 3.940 0.960 ;
        RECT  3.140 2.230 3.865 2.390 ;
        RECT  2.965 0.800 3.730 0.960 ;
        RECT  3.490 1.580 3.650 1.880 ;
        RECT  2.540 1.720 3.490 1.880 ;
        RECT  3.190 0.310 3.450 0.620 ;
        RECT  2.980 2.230 3.140 2.560 ;
        RECT  2.965 1.280 3.100 1.540 ;
        RECT  0.680 2.400 2.980 2.560 ;
        RECT  2.805 0.410 2.965 1.540 ;
        RECT  2.730 0.410 2.805 0.670 ;
        RECT  1.625 1.310 2.805 1.470 ;
        RECT  1.110 2.060 2.800 2.220 ;
        RECT  2.280 1.685 2.540 1.880 ;
        RECT  1.445 0.460 2.430 0.620 ;
        RECT  1.445 1.685 2.280 1.845 ;
        RECT  1.285 0.460 1.445 1.845 ;
        RECT  0.940 0.460 1.285 0.620 ;
        RECT  1.160 1.585 1.285 1.845 ;
        RECT  0.975 2.030 1.110 2.220 ;
        RECT  0.975 0.800 1.090 1.060 ;
        RECT  0.815 0.800 0.975 2.220 ;
        RECT  0.680 0.310 0.940 0.620 ;
    END
END DFFSX4MTH

MACRO DFFTRX1MTH
    CLASS CORE ;
    FOREIGN DFFTRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.585 1.170 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.785 0.815 7.845 0.975 ;
        RECT  7.525 0.815 7.785 2.245 ;
        RECT  7.480 1.290 7.525 1.580 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 1.290 8.920 1.580 ;
        RECT  8.635 0.745 8.895 2.255 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.780 1.290 1.130 1.695 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.525 1.295 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.345 -0.130 9.020 0.130 ;
        RECT  7.745 -0.130 8.345 0.280 ;
        RECT  6.765 -0.130 7.745 0.130 ;
        RECT  6.505 -0.130 6.765 0.300 ;
        RECT  4.875 -0.130 6.505 0.130 ;
        RECT  4.615 -0.130 4.875 0.685 ;
        RECT  2.785 -0.130 4.615 0.130 ;
        RECT  2.525 -0.130 2.785 0.335 ;
        RECT  0.385 -0.130 2.525 0.130 ;
        RECT  0.125 -0.130 0.385 0.700 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.340 2.740 9.020 3.000 ;
        RECT  8.080 1.835 8.340 3.000 ;
        RECT  6.705 2.740 8.080 3.000 ;
        RECT  6.445 2.515 6.705 3.000 ;
        RECT  4.485 2.740 6.445 3.000 ;
        RECT  4.225 2.050 4.485 3.000 ;
        RECT  1.235 2.740 4.225 3.000 ;
        RECT  0.635 2.380 1.235 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.285 0.475 8.445 1.610 ;
        RECT  7.295 0.475 8.285 0.635 ;
        RECT  7.135 0.475 7.295 2.295 ;
        RECT  7.105 0.475 7.135 0.755 ;
        RECT  6.685 1.455 7.135 1.615 ;
        RECT  7.015 2.035 7.135 2.295 ;
        RECT  6.795 0.875 6.955 1.135 ;
        RECT  6.345 0.875 6.795 1.035 ;
        RECT  6.525 1.355 6.685 1.615 ;
        RECT  6.185 0.875 6.345 2.195 ;
        RECT  5.945 0.875 6.185 1.035 ;
        RECT  5.915 2.035 6.185 2.195 ;
        RECT  5.845 1.465 6.005 1.725 ;
        RECT  5.785 0.495 5.945 1.035 ;
        RECT  5.755 2.035 5.915 2.295 ;
        RECT  5.575 1.565 5.845 1.725 ;
        RECT  5.415 1.565 5.575 2.405 ;
        RECT  4.855 2.245 5.415 2.405 ;
        RECT  5.235 0.655 5.375 1.025 ;
        RECT  5.215 0.655 5.235 2.065 ;
        RECT  5.075 0.865 5.215 2.065 ;
        RECT  4.605 0.865 5.075 1.025 ;
        RECT  4.695 1.345 4.855 2.405 ;
        RECT  4.265 1.345 4.695 1.505 ;
        RECT  4.445 0.865 4.605 1.165 ;
        RECT  3.925 1.700 4.515 1.860 ;
        RECT  4.105 0.310 4.265 1.505 ;
        RECT  3.365 0.310 4.105 0.470 ;
        RECT  3.765 0.650 3.925 2.455 ;
        RECT  3.665 0.650 3.765 0.810 ;
        RECT  3.055 2.295 3.765 2.455 ;
        RECT  3.365 1.055 3.505 1.315 ;
        RECT  3.205 0.310 3.365 2.085 ;
        RECT  3.145 0.490 3.205 0.750 ;
        RECT  3.155 1.695 3.205 2.085 ;
        RECT  2.285 1.925 3.155 2.085 ;
        RECT  2.895 2.295 3.055 2.560 ;
        RECT  2.865 0.955 3.025 1.215 ;
        RECT  1.845 2.400 2.895 2.560 ;
        RECT  2.705 0.540 2.865 1.650 ;
        RECT  1.865 0.540 2.705 0.700 ;
        RECT  2.165 1.490 2.705 1.650 ;
        RECT  2.025 1.925 2.285 2.220 ;
        RECT  1.705 0.540 1.865 1.185 ;
        RECT  1.685 1.515 1.845 2.560 ;
        RECT  1.525 1.515 1.685 1.675 ;
        RECT  1.365 0.440 1.525 1.675 ;
        RECT  0.385 1.875 1.325 2.035 ;
        RECT  0.225 1.875 0.385 2.500 ;
        RECT  0.125 2.340 0.225 2.500 ;
    END
END DFFTRX1MTH

MACRO DFFTRX2MTH
    CLASS CORE ;
    FOREIGN DFFTRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.585 1.170 ;
        END
        AntennaGateArea 0.0637 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.740 0.815 7.815 0.975 ;
        RECT  7.740 1.685 7.785 2.285 ;
        RECT  7.480 0.815 7.740 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 1.290 8.920 1.580 ;
        RECT  8.635 0.425 8.895 2.425 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.780 1.290 1.130 1.695 ;
        END
        AntennaGateArea 0.0676 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 0.880 2.485 1.295 ;
        END
        AntennaGateArea 0.1014 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 -0.130 9.020 0.130 ;
        RECT  8.095 -0.130 8.355 0.250 ;
        RECT  6.715 -0.130 8.095 0.130 ;
        RECT  6.455 -0.130 6.715 0.300 ;
        RECT  4.885 -0.130 6.455 0.130 ;
        RECT  4.625 -0.130 4.885 0.685 ;
        RECT  2.735 -0.130 4.625 0.130 ;
        RECT  2.475 -0.130 2.735 0.300 ;
        RECT  0.385 -0.130 2.475 0.130 ;
        RECT  0.125 -0.130 0.385 0.700 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.340 2.740 9.020 3.000 ;
        RECT  8.080 1.835 8.340 3.000 ;
        RECT  6.705 2.740 8.080 3.000 ;
        RECT  6.445 2.515 6.705 3.000 ;
        RECT  4.485 2.740 6.445 3.000 ;
        RECT  4.225 2.050 4.485 3.000 ;
        RECT  1.235 2.740 4.225 3.000 ;
        RECT  0.635 2.380 1.235 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.295 0.475 8.455 1.545 ;
        RECT  7.275 0.475 8.295 0.635 ;
        RECT  7.115 0.475 7.275 2.295 ;
        RECT  7.085 0.475 7.115 0.755 ;
        RECT  6.685 1.455 7.115 1.615 ;
        RECT  7.015 2.035 7.115 2.295 ;
        RECT  6.755 0.875 6.915 1.135 ;
        RECT  6.345 0.875 6.755 1.035 ;
        RECT  6.525 1.355 6.685 1.615 ;
        RECT  6.185 0.875 6.345 2.195 ;
        RECT  5.915 0.875 6.185 1.035 ;
        RECT  5.915 2.035 6.185 2.195 ;
        RECT  5.845 1.595 6.005 1.855 ;
        RECT  5.755 0.525 5.915 1.035 ;
        RECT  5.755 2.035 5.915 2.295 ;
        RECT  5.575 1.695 5.845 1.855 ;
        RECT  5.415 1.695 5.575 2.405 ;
        RECT  4.855 2.245 5.415 2.405 ;
        RECT  5.245 0.625 5.405 1.025 ;
        RECT  5.235 0.865 5.245 1.025 ;
        RECT  5.075 0.865 5.235 2.065 ;
        RECT  4.585 0.865 5.075 1.025 ;
        RECT  4.695 1.345 4.855 2.405 ;
        RECT  4.225 1.345 4.695 1.505 ;
        RECT  4.425 0.865 4.585 1.165 ;
        RECT  3.885 1.700 4.515 1.860 ;
        RECT  4.065 0.310 4.225 1.505 ;
        RECT  3.365 0.310 4.065 0.470 ;
        RECT  3.725 0.650 3.885 2.455 ;
        RECT  3.615 0.650 3.725 0.810 ;
        RECT  3.015 2.295 3.725 2.455 ;
        RECT  3.365 1.055 3.505 1.315 ;
        RECT  3.205 0.310 3.365 2.085 ;
        RECT  3.095 0.450 3.205 0.710 ;
        RECT  3.115 1.695 3.205 2.085 ;
        RECT  2.285 1.925 3.115 2.085 ;
        RECT  2.865 0.955 3.025 1.215 ;
        RECT  2.855 2.295 3.015 2.560 ;
        RECT  2.705 0.490 2.865 1.650 ;
        RECT  1.845 2.400 2.855 2.560 ;
        RECT  1.930 0.490 2.705 0.650 ;
        RECT  2.165 1.490 2.705 1.650 ;
        RECT  2.025 1.925 2.285 2.220 ;
        RECT  1.770 0.490 1.930 1.200 ;
        RECT  1.685 1.515 1.845 2.560 ;
        RECT  1.525 1.515 1.685 1.675 ;
        RECT  1.365 0.440 1.525 1.675 ;
        RECT  0.385 1.875 1.325 2.035 ;
        RECT  0.225 1.875 0.385 2.500 ;
        RECT  0.125 2.340 0.225 2.500 ;
    END
END DFFTRX2MTH

MACRO DFFTRX4MTH
    CLASS CORE ;
    FOREIGN DFFTRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 0.915 1.170 1.135 ;
        RECT  0.445 0.975 0.470 1.135 ;
        END
        AntennaGateArea 0.0975 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.325 0.815 10.585 2.415 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 1.290 11.790 1.580 ;
        RECT  11.405 0.420 11.665 2.425 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.670 1.330 1.245 1.665 ;
        END
        AntennaGateArea 0.1313 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 0.880 2.770 1.295 ;
        END
        AntennaGateArea 0.1521 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 -0.130 12.300 0.130 ;
        RECT  11.915 -0.130 12.175 1.020 ;
        RECT  11.125 -0.130 11.915 0.130 ;
        RECT  10.865 -0.130 11.125 0.285 ;
        RECT  10.045 -0.130 10.865 0.130 ;
        RECT  9.785 -0.130 10.045 0.250 ;
        RECT  9.045 -0.130 9.785 0.130 ;
        RECT  8.445 -0.130 9.045 0.250 ;
        RECT  6.460 -0.130 8.445 0.130 ;
        RECT  6.300 -0.130 6.460 1.035 ;
        RECT  5.100 -0.130 6.300 0.130 ;
        RECT  4.840 -0.130 5.100 0.575 ;
        RECT  3.095 -0.130 4.840 0.130 ;
        RECT  2.495 -0.130 3.095 0.300 ;
        RECT  0.535 -0.130 2.495 0.130 ;
        RECT  0.275 -0.130 0.535 0.575 ;
        RECT  0.000 -0.130 0.275 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 2.740 12.300 3.000 ;
        RECT  11.915 1.825 12.175 3.000 ;
        RECT  11.125 2.740 11.915 3.000 ;
        RECT  10.865 1.825 11.125 3.000 ;
        RECT  10.075 2.740 10.865 3.000 ;
        RECT  9.815 1.825 10.075 3.000 ;
        RECT  9.055 2.740 9.815 3.000 ;
        RECT  8.795 1.890 9.055 3.000 ;
        RECT  6.570 2.740 8.795 3.000 ;
        RECT  6.410 1.955 6.570 3.000 ;
        RECT  5.550 2.740 6.410 3.000 ;
        RECT  5.390 1.955 5.550 3.000 ;
        RECT  4.500 2.740 5.390 3.000 ;
        RECT  4.340 2.025 4.500 3.000 ;
        RECT  2.965 2.740 4.340 3.000 ;
        RECT  2.365 2.620 2.965 3.000 ;
        RECT  1.635 2.740 2.365 3.000 ;
        RECT  0.695 2.620 1.635 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.065 0.475 11.225 1.575 ;
        RECT  9.925 0.475 11.065 0.635 ;
        RECT  9.765 0.475 9.925 0.965 ;
        RECT  9.515 0.805 9.765 0.965 ;
        RECT  9.515 1.890 9.565 2.150 ;
        RECT  9.355 0.805 9.515 2.150 ;
        RECT  9.190 0.395 9.450 0.590 ;
        RECT  8.920 1.135 9.355 1.295 ;
        RECT  9.305 1.890 9.355 2.150 ;
        RECT  8.580 0.430 9.190 0.590 ;
        RECT  8.760 1.135 8.920 1.395 ;
        RECT  8.420 0.430 8.580 2.065 ;
        RECT  8.040 0.430 8.420 0.590 ;
        RECT  8.110 1.905 8.420 2.065 ;
        RECT  8.080 1.095 8.240 1.725 ;
        RECT  7.950 1.905 8.110 2.505 ;
        RECT  7.480 1.095 8.080 1.255 ;
        RECT  7.780 0.430 8.040 0.690 ;
        RECT  7.080 2.345 7.950 2.505 ;
        RECT  7.430 1.555 7.590 2.090 ;
        RECT  7.320 0.565 7.480 1.255 ;
        RECT  7.140 1.555 7.430 1.715 ;
        RECT  6.800 0.565 7.320 0.725 ;
        RECT  6.980 0.905 7.140 1.715 ;
        RECT  6.920 1.905 7.080 2.505 ;
        RECT  6.060 1.555 6.980 1.715 ;
        RECT  6.640 0.565 6.800 1.375 ;
        RECT  6.120 1.215 6.640 1.375 ;
        RECT  5.960 0.565 6.120 1.375 ;
        RECT  5.900 1.555 6.060 2.180 ;
        RECT  5.440 0.565 5.960 0.725 ;
        RECT  5.780 1.555 5.900 1.715 ;
        RECT  5.620 0.905 5.780 1.715 ;
        RECT  5.040 1.095 5.620 1.255 ;
        RECT  5.280 0.565 5.440 0.915 ;
        RECT  4.490 0.755 5.280 0.915 ;
        RECT  4.880 1.095 5.040 2.180 ;
        RECT  4.640 1.095 4.880 1.255 ;
        RECT  4.140 1.575 4.660 1.735 ;
        RECT  4.330 0.310 4.490 0.915 ;
        RECT  3.485 0.310 4.330 0.470 ;
        RECT  3.980 0.650 4.140 2.440 ;
        RECT  1.815 2.280 3.980 2.440 ;
        RECT  3.485 0.920 3.800 1.080 ;
        RECT  3.455 0.310 3.485 1.080 ;
        RECT  3.325 0.310 3.455 2.100 ;
        RECT  3.295 0.920 3.325 2.100 ;
        RECT  1.995 1.940 3.295 2.100 ;
        RECT  2.955 0.540 3.115 1.730 ;
        RECT  2.025 0.540 2.955 0.700 ;
        RECT  2.255 1.570 2.955 1.730 ;
        RECT  1.865 0.540 2.025 1.185 ;
        RECT  1.685 1.890 1.815 2.440 ;
        RECT  1.525 0.465 1.685 2.440 ;
        RECT  1.405 0.465 1.525 0.725 ;
        RECT  1.145 1.875 1.305 2.135 ;
        RECT  0.525 1.975 1.145 2.135 ;
        RECT  0.365 1.975 0.525 2.485 ;
        RECT  0.185 2.325 0.365 2.485 ;
    END
END DFFTRX4MTH

MACRO DFFX1MTH
    CLASS CORE ;
    FOREIGN DFFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 0.735 6.565 1.170 ;
        RECT  6.095 1.930 6.565 2.090 ;
        RECT  6.095 1.010 6.250 1.170 ;
        RECT  5.935 1.010 6.095 2.090 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 1.290 8.100 1.580 ;
        RECT  7.865 0.755 8.075 2.195 ;
        RECT  7.815 0.755 7.865 1.015 ;
        RECT  7.815 1.935 7.865 2.195 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.090 0.400 1.675 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.000 1.715 2.400 2.065 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.525 -0.130 8.200 0.130 ;
        RECT  6.925 -0.130 7.525 0.365 ;
        RECT  6.495 -0.130 6.925 0.130 ;
        RECT  5.895 -0.130 6.495 0.385 ;
        RECT  4.385 -0.130 5.895 0.130 ;
        RECT  4.125 -0.130 4.385 0.345 ;
        RECT  0.730 -0.130 4.125 0.130 ;
        RECT  0.130 -0.130 0.730 0.350 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 2.740 8.200 3.000 ;
        RECT  6.935 2.620 7.535 3.000 ;
        RECT  6.495 2.740 6.935 3.000 ;
        RECT  5.895 2.620 6.495 3.000 ;
        RECT  1.960 2.740 5.895 3.000 ;
        RECT  1.700 2.620 1.960 3.000 ;
        RECT  0.385 2.740 1.700 3.000 ;
        RECT  0.125 2.510 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.460 1.380 7.560 1.640 ;
        RECT  7.300 1.380 7.460 2.430 ;
        RECT  5.755 2.270 7.300 2.430 ;
        RECT  6.915 0.760 7.075 2.035 ;
        RECT  6.815 0.760 6.915 1.020 ;
        RECT  6.815 1.535 6.915 2.035 ;
        RECT  6.535 1.535 6.815 1.695 ;
        RECT  6.375 1.350 6.535 1.695 ;
        RECT  6.275 1.350 6.375 1.510 ;
        RECT  5.595 0.680 5.755 2.430 ;
        RECT  5.005 0.680 5.595 0.840 ;
        RECT  5.005 2.200 5.595 2.430 ;
        RECT  5.255 1.020 5.415 1.280 ;
        RECT  5.070 1.120 5.255 1.280 ;
        RECT  4.910 1.120 5.070 2.020 ;
        RECT  4.730 0.310 5.065 0.470 ;
        RECT  4.675 1.860 4.910 2.020 ;
        RECT  4.570 0.310 4.730 1.155 ;
        RECT  4.515 1.860 4.675 2.545 ;
        RECT  4.335 1.335 4.585 1.495 ;
        RECT  3.905 0.995 4.570 1.155 ;
        RECT  2.540 2.385 4.515 2.545 ;
        RECT  4.175 1.335 4.335 2.205 ;
        RECT  2.960 2.045 4.175 2.205 ;
        RECT  3.905 1.705 3.935 1.865 ;
        RECT  3.745 0.310 3.905 1.865 ;
        RECT  1.240 0.310 3.745 0.470 ;
        RECT  3.675 1.705 3.745 1.865 ;
        RECT  3.285 0.665 3.445 1.535 ;
        RECT  3.185 0.665 3.285 0.825 ;
        RECT  2.960 1.375 3.285 1.535 ;
        RECT  1.080 1.035 3.105 1.195 ;
        RECT  2.800 1.375 2.960 2.205 ;
        RECT  1.550 1.375 2.800 1.535 ;
        RECT  2.750 2.045 2.800 2.205 ;
        RECT  2.380 2.280 2.540 2.545 ;
        RECT  0.950 0.650 2.460 0.810 ;
        RECT  1.420 2.280 2.380 2.440 ;
        RECT  1.260 2.280 1.420 2.535 ;
        RECT  1.070 2.350 1.260 2.535 ;
        RECT  0.920 0.990 1.080 2.170 ;
        RECT  0.740 2.350 1.070 2.510 ;
        RECT  0.740 0.530 0.950 0.810 ;
        RECT  0.670 0.530 0.740 2.510 ;
        RECT  0.580 0.650 0.670 2.510 ;
    END
END DFFX1MTH

MACRO DFFX2MTH
    CLASS CORE ;
    FOREIGN DFFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.485 1.290 8.510 1.580 ;
        RECT  8.225 0.400 8.485 2.355 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.580 1.685 7.690 1.990 ;
        RECT  7.370 0.765 7.580 1.990 ;
        RECT  7.275 0.765 7.370 1.025 ;
        RECT  7.245 1.685 7.370 1.990 ;
        END
        AntennaDiffArea 0.478 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.100 0.395 1.655 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.740 2.470 1.950 ;
        END
        AntennaGateArea 0.0871 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 -0.130 8.610 0.130 ;
        RECT  7.685 -0.130 7.945 0.515 ;
        RECT  6.915 -0.130 7.685 0.130 ;
        RECT  6.315 -0.130 6.915 0.250 ;
        RECT  4.575 -0.130 6.315 0.130 ;
        RECT  4.315 -0.130 4.575 0.650 ;
        RECT  0.725 -0.130 4.315 0.130 ;
        RECT  0.125 -0.130 0.725 0.350 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 2.740 8.610 3.000 ;
        RECT  7.685 2.550 7.945 3.000 ;
        RECT  6.965 2.740 7.685 3.000 ;
        RECT  6.365 2.510 6.965 3.000 ;
        RECT  4.765 2.740 6.365 3.000 ;
        RECT  4.165 2.620 4.765 3.000 ;
        RECT  3.985 2.740 4.165 3.000 ;
        RECT  3.385 2.620 3.985 3.000 ;
        RECT  2.100 2.740 3.385 3.000 ;
        RECT  1.840 2.620 2.100 3.000 ;
        RECT  0.460 2.740 1.840 3.000 ;
        RECT  0.200 1.990 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.875 1.270 8.035 2.330 ;
        RECT  6.335 2.170 7.875 2.330 ;
        RECT  7.070 1.200 7.120 1.460 ;
        RECT  6.910 0.430 7.070 1.460 ;
        RECT  5.995 0.430 6.910 0.590 ;
        RECT  6.860 1.200 6.910 1.460 ;
        RECT  6.335 0.815 6.495 0.975 ;
        RECT  6.335 1.685 6.485 1.945 ;
        RECT  6.175 0.815 6.335 2.330 ;
        RECT  5.835 0.430 5.995 2.235 ;
        RECT  5.345 0.430 5.835 0.590 ;
        RECT  5.595 2.075 5.835 2.235 ;
        RECT  5.495 0.880 5.655 1.385 ;
        RECT  5.435 2.075 5.595 2.395 ;
        RECT  5.445 1.220 5.495 1.385 ;
        RECT  5.255 1.220 5.445 1.880 ;
        RECT  5.185 0.430 5.345 0.700 ;
        RECT  5.095 1.220 5.255 2.440 ;
        RECT  3.940 0.880 5.225 1.040 ;
        RECT  4.120 1.220 5.095 1.380 ;
        RECT  1.605 2.280 5.095 2.440 ;
        RECT  4.755 1.670 4.915 2.100 ;
        RECT  3.085 1.940 4.755 2.100 ;
        RECT  3.940 1.600 4.545 1.760 ;
        RECT  3.780 0.310 3.940 1.760 ;
        RECT  1.285 0.310 3.780 0.470 ;
        RECT  3.385 0.650 3.545 1.545 ;
        RECT  3.220 0.650 3.385 0.810 ;
        RECT  3.085 1.385 3.385 1.545 ;
        RECT  1.260 1.035 3.205 1.195 ;
        RECT  2.925 1.385 3.085 2.100 ;
        RECT  1.730 1.385 2.925 1.545 ;
        RECT  0.975 0.650 2.500 0.810 ;
        RECT  1.445 2.280 1.605 2.545 ;
        RECT  0.920 2.385 1.445 2.545 ;
        RECT  1.175 1.035 1.260 2.165 ;
        RECT  1.100 0.990 1.175 2.165 ;
        RECT  0.915 0.990 1.100 1.195 ;
        RECT  0.735 0.555 0.975 0.810 ;
        RECT  0.760 1.545 0.920 2.545 ;
        RECT  0.735 1.545 0.760 1.705 ;
        RECT  0.685 0.555 0.735 1.705 ;
        RECT  0.575 0.650 0.685 1.705 ;
    END
END DFFX2MTH

MACRO DFFX4MTH
    CLASS CORE ;
    FOREIGN DFFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.745 1.290 8.920 1.580 ;
        RECT  8.485 0.400 8.745 2.355 ;
        END
        AntennaDiffArea 0.68 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.420 0.425 7.690 1.900 ;
        RECT  7.360 1.740 7.420 1.900 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.150 0.395 1.700 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.740 2.470 1.960 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.295 -0.130 9.430 0.130 ;
        RECT  9.035 -0.130 9.295 1.025 ;
        RECT  8.195 -0.130 9.035 0.130 ;
        RECT  7.935 -0.130 8.195 0.985 ;
        RECT  7.125 -0.130 7.935 0.130 ;
        RECT  6.185 -0.130 7.125 0.250 ;
        RECT  4.565 -0.130 6.185 0.130 ;
        RECT  4.305 -0.130 4.565 0.535 ;
        RECT  1.090 -0.130 4.305 0.130 ;
        RECT  0.150 -0.130 1.090 0.310 ;
        RECT  0.000 -0.130 0.150 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.295 2.740 9.430 3.000 ;
        RECT  9.035 1.885 9.295 3.000 ;
        RECT  8.165 2.740 9.035 3.000 ;
        RECT  7.905 2.420 8.165 3.000 ;
        RECT  6.970 2.740 7.905 3.000 ;
        RECT  6.370 2.445 6.970 3.000 ;
        RECT  2.100 2.740 6.370 3.000 ;
        RECT  1.840 2.620 2.100 3.000 ;
        RECT  0.410 2.740 1.840 3.000 ;
        RECT  0.150 1.890 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.145 1.235 8.305 2.240 ;
        RECT  6.550 2.080 8.145 2.240 ;
        RECT  7.175 1.230 7.225 1.490 ;
        RECT  7.015 0.435 7.175 1.490 ;
        RECT  6.040 0.435 7.015 0.595 ;
        RECT  6.965 1.230 7.015 1.490 ;
        RECT  6.550 0.815 6.715 0.975 ;
        RECT  6.390 0.815 6.550 2.240 ;
        RECT  6.315 0.815 6.390 0.975 ;
        RECT  6.370 1.310 6.390 2.240 ;
        RECT  6.220 1.310 6.370 1.570 ;
        RECT  5.880 0.370 6.040 2.235 ;
        RECT  5.215 0.370 5.880 0.530 ;
        RECT  5.605 2.075 5.880 2.235 ;
        RECT  5.515 0.715 5.675 1.715 ;
        RECT  5.445 2.075 5.605 2.385 ;
        RECT  4.230 0.715 5.515 0.875 ;
        RECT  5.260 1.555 5.515 1.715 ;
        RECT  5.100 1.555 5.260 2.545 ;
        RECT  4.570 1.075 5.245 1.235 ;
        RECT  2.640 2.385 5.100 2.545 ;
        RECT  4.760 1.505 4.920 2.205 ;
        RECT  3.235 2.045 4.760 2.205 ;
        RECT  4.410 1.075 4.570 1.865 ;
        RECT  3.890 1.705 4.410 1.865 ;
        RECT  4.070 0.715 4.230 1.365 ;
        RECT  3.890 0.325 3.990 0.545 ;
        RECT  3.730 0.325 3.890 1.865 ;
        RECT  1.290 0.325 3.730 0.485 ;
        RECT  3.380 0.665 3.540 1.550 ;
        RECT  3.220 0.665 3.380 0.825 ;
        RECT  3.235 1.390 3.380 1.550 ;
        RECT  3.075 1.390 3.235 2.205 ;
        RECT  2.935 1.015 3.195 1.210 ;
        RECT  1.730 1.390 3.075 1.550 ;
        RECT  1.260 1.015 2.935 1.175 ;
        RECT  2.380 2.265 2.640 2.545 ;
        RECT  0.950 0.665 2.500 0.825 ;
        RECT  1.605 2.265 2.380 2.425 ;
        RECT  1.445 2.265 1.605 2.470 ;
        RECT  0.870 2.310 1.445 2.470 ;
        RECT  1.260 1.940 1.310 2.100 ;
        RECT  1.100 1.015 1.260 2.100 ;
        RECT  0.920 1.015 1.100 1.195 ;
        RECT  1.050 1.940 1.100 2.100 ;
        RECT  0.740 0.490 0.950 0.825 ;
        RECT  0.740 1.545 0.870 2.470 ;
        RECT  0.710 0.490 0.740 2.470 ;
        RECT  0.690 0.490 0.710 1.705 ;
        RECT  0.580 0.665 0.690 1.705 ;
    END
END DFFX4MTH

MACRO DLY1X1MTH
    CLASS CORE ;
    FOREIGN DLY1X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.765 3.180 2.380 ;
        RECT  2.895 0.765 2.970 1.025 ;
        RECT  2.895 2.120 2.970 2.380 ;
        END
        AntennaDiffArea 0.279 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.150 0.815 1.610 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.075 -0.130 3.280 0.130 ;
        RECT  2.475 -0.130 3.075 0.450 ;
        RECT  1.265 -0.130 2.475 0.130 ;
        RECT  0.325 -0.130 1.265 0.460 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 2.740 3.280 3.000 ;
        RECT  0.325 2.300 1.265 3.000 ;
        RECT  0.000 2.740 0.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.710 1.225 2.790 1.485 ;
        RECT  2.550 0.655 2.710 2.460 ;
        RECT  2.155 0.655 2.550 0.815 ;
        RECT  1.775 2.300 2.550 2.460 ;
        RECT  1.775 1.035 2.270 1.535 ;
        RECT  1.995 0.420 2.155 0.815 ;
        RECT  1.775 0.420 1.995 0.580 ;
        RECT  1.515 0.320 1.775 0.580 ;
        RECT  1.515 0.830 1.775 2.015 ;
        RECT  1.515 2.300 1.775 2.560 ;
        RECT  1.035 1.130 1.295 1.950 ;
        RECT  0.385 1.790 1.035 1.950 ;
        RECT  0.285 0.710 0.385 0.970 ;
        RECT  0.285 1.790 0.385 2.050 ;
        RECT  0.125 0.710 0.285 2.050 ;
    END
END DLY1X1MTH

MACRO DLY1X4MTH
    CLASS CORE ;
    FOREIGN DLY1X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.930 1.045 4.000 1.730 ;
        RECT  3.670 0.610 3.930 1.730 ;
        RECT  3.455 1.570 3.670 1.730 ;
        RECT  3.195 1.570 3.455 2.435 ;
        END
        AntennaDiffArea 0.551 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 0.920 0.760 1.580 ;
        END
        AntennaGateArea 0.13 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 -0.130 4.100 0.130 ;
        RECT  3.100 -0.130 3.360 0.725 ;
        RECT  0.905 -0.130 3.100 0.130 ;
        RECT  0.645 -0.130 0.905 0.740 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 1.910 3.975 3.000 ;
        RECT  1.125 2.740 3.715 3.000 ;
        RECT  0.185 2.535 1.125 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.005 1.230 3.450 1.390 ;
        RECT  2.845 0.905 3.005 2.355 ;
        RECT  2.315 0.905 2.845 1.065 ;
        RECT  2.115 2.195 2.845 2.355 ;
        RECT  2.300 1.245 2.560 1.745 ;
        RECT  2.055 0.765 2.315 1.065 ;
        RECT  1.755 1.245 2.300 1.495 ;
        RECT  1.855 2.195 2.115 2.455 ;
        RECT  1.755 0.455 1.805 0.715 ;
        RECT  1.505 0.455 1.755 1.945 ;
        RECT  1.455 1.685 1.505 1.945 ;
        RECT  1.190 1.025 1.290 1.525 ;
        RECT  1.030 1.025 1.190 1.925 ;
        RECT  0.385 1.765 1.030 1.925 ;
        RECT  0.285 0.480 0.385 0.740 ;
        RECT  0.285 1.765 0.385 2.085 ;
        RECT  0.125 0.480 0.285 2.085 ;
    END
END DLY1X4MTH

MACRO DLY2X1MTH
    CLASS CORE ;
    FOREIGN DLY2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.765 3.180 2.380 ;
        RECT  2.895 0.765 2.970 1.025 ;
        RECT  2.895 2.120 2.970 2.380 ;
        END
        AntennaDiffArea 0.275 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.150 0.815 1.610 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.075 -0.130 3.280 0.130 ;
        RECT  2.475 -0.130 3.075 0.450 ;
        RECT  1.265 -0.130 2.475 0.130 ;
        RECT  0.325 -0.130 1.265 0.460 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 2.740 3.280 3.000 ;
        RECT  0.325 2.300 1.265 3.000 ;
        RECT  0.000 2.740 0.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.710 1.225 2.790 1.485 ;
        RECT  2.550 0.655 2.710 2.460 ;
        RECT  2.155 0.655 2.550 0.815 ;
        RECT  1.775 2.300 2.550 2.460 ;
        RECT  1.775 1.035 2.270 1.535 ;
        RECT  1.995 0.420 2.155 0.815 ;
        RECT  1.775 0.420 1.995 0.580 ;
        RECT  1.515 0.320 1.775 0.580 ;
        RECT  1.515 0.830 1.775 2.015 ;
        RECT  1.515 2.300 1.775 2.560 ;
        RECT  1.035 1.130 1.315 1.950 ;
        RECT  0.385 1.790 1.035 1.950 ;
        RECT  0.285 0.710 0.385 0.970 ;
        RECT  0.285 1.790 0.385 2.050 ;
        RECT  0.125 0.710 0.285 2.050 ;
    END
END DLY2X1MTH

MACRO DLY2X4MTH
    CLASS CORE ;
    FOREIGN DLY2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.930 1.045 4.000 1.730 ;
        RECT  3.670 0.610 3.930 1.730 ;
        RECT  3.455 1.570 3.670 1.730 ;
        RECT  3.195 1.570 3.455 2.435 ;
        END
        AntennaDiffArea 0.555 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 0.920 0.760 1.580 ;
        END
        AntennaGateArea 0.13 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 -0.130 4.100 0.130 ;
        RECT  3.100 -0.130 3.360 0.725 ;
        RECT  0.905 -0.130 3.100 0.130 ;
        RECT  0.645 -0.130 0.905 0.740 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 1.915 3.975 3.000 ;
        RECT  1.130 2.740 3.715 3.000 ;
        RECT  0.190 2.535 1.130 3.000 ;
        RECT  0.000 2.740 0.190 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.005 1.230 3.450 1.390 ;
        RECT  2.845 0.905 3.005 2.355 ;
        RECT  2.315 0.905 2.845 1.065 ;
        RECT  2.115 2.195 2.845 2.355 ;
        RECT  2.300 1.245 2.560 1.745 ;
        RECT  2.055 0.765 2.315 1.065 ;
        RECT  1.755 1.245 2.300 1.495 ;
        RECT  1.855 2.195 2.115 2.455 ;
        RECT  1.755 0.455 1.805 0.715 ;
        RECT  1.505 0.455 1.755 1.945 ;
        RECT  1.455 1.685 1.505 1.945 ;
        RECT  1.190 1.025 1.290 1.525 ;
        RECT  1.030 1.025 1.190 1.925 ;
        RECT  0.385 1.765 1.030 1.925 ;
        RECT  0.285 0.480 0.385 0.740 ;
        RECT  0.285 1.765 0.385 2.085 ;
        RECT  0.125 0.480 0.285 2.085 ;
    END
END DLY2X4MTH

MACRO DLY3X1MTH
    CLASS CORE ;
    FOREIGN DLY3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.765 3.180 2.380 ;
        RECT  2.895 0.765 2.970 1.025 ;
        RECT  2.895 2.120 2.970 2.380 ;
        END
        AntennaDiffArea 0.275 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.150 0.815 1.610 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.075 -0.130 3.280 0.130 ;
        RECT  2.475 -0.130 3.075 0.450 ;
        RECT  1.265 -0.130 2.475 0.130 ;
        RECT  0.325 -0.130 1.265 0.460 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 2.740 3.280 3.000 ;
        RECT  0.325 2.300 1.265 3.000 ;
        RECT  0.000 2.740 0.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.710 1.225 2.790 1.485 ;
        RECT  2.550 0.655 2.710 2.460 ;
        RECT  2.155 0.655 2.550 0.815 ;
        RECT  1.775 2.300 2.550 2.460 ;
        RECT  1.775 1.035 2.270 1.535 ;
        RECT  1.995 0.420 2.155 0.815 ;
        RECT  1.775 0.420 1.995 0.580 ;
        RECT  1.515 0.320 1.775 0.580 ;
        RECT  1.515 0.830 1.775 2.015 ;
        RECT  1.515 2.300 1.775 2.560 ;
        RECT  1.035 1.130 1.315 1.950 ;
        RECT  0.385 1.790 1.035 1.950 ;
        RECT  0.285 0.710 0.385 0.970 ;
        RECT  0.285 1.790 0.385 2.050 ;
        RECT  0.125 0.710 0.285 2.050 ;
    END
END DLY3X1MTH

MACRO DLY3X4MTH
    CLASS CORE ;
    FOREIGN DLY3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.930 1.045 4.000 1.730 ;
        RECT  3.670 0.610 3.930 1.730 ;
        RECT  3.455 1.570 3.670 1.730 ;
        RECT  3.195 1.570 3.455 2.435 ;
        END
        AntennaDiffArea 0.555 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 0.920 0.760 1.580 ;
        END
        AntennaGateArea 0.13 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 -0.130 4.100 0.130 ;
        RECT  3.100 -0.130 3.360 0.725 ;
        RECT  0.905 -0.130 3.100 0.130 ;
        RECT  0.645 -0.130 0.905 0.740 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 1.915 3.975 3.000 ;
        RECT  1.125 2.740 3.715 3.000 ;
        RECT  0.185 2.535 1.125 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.005 1.230 3.450 1.390 ;
        RECT  2.845 0.905 3.005 2.355 ;
        RECT  2.315 0.905 2.845 1.065 ;
        RECT  2.115 2.195 2.845 2.355 ;
        RECT  2.300 1.245 2.560 1.745 ;
        RECT  2.055 0.765 2.315 1.065 ;
        RECT  1.755 1.245 2.300 1.495 ;
        RECT  1.855 2.195 2.115 2.455 ;
        RECT  1.755 0.455 1.805 0.715 ;
        RECT  1.505 0.455 1.755 1.945 ;
        RECT  1.455 1.685 1.505 1.945 ;
        RECT  1.190 1.025 1.290 1.525 ;
        RECT  1.030 1.025 1.190 1.925 ;
        RECT  0.385 1.765 1.030 1.925 ;
        RECT  0.285 0.480 0.385 0.740 ;
        RECT  0.285 1.765 0.385 2.085 ;
        RECT  0.125 0.480 0.285 2.085 ;
    END
END DLY3X4MTH

MACRO DLY4X1MTH
    CLASS CORE ;
    FOREIGN DLY4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.765 3.180 2.380 ;
        RECT  2.895 0.765 2.970 1.025 ;
        RECT  2.895 2.120 2.970 2.380 ;
        END
        AntennaDiffArea 0.279 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.150 0.815 1.610 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.075 -0.130 3.280 0.130 ;
        RECT  2.475 -0.130 3.075 0.450 ;
        RECT  1.265 -0.130 2.475 0.130 ;
        RECT  0.325 -0.130 1.265 0.460 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 2.740 3.280 3.000 ;
        RECT  0.325 2.300 1.265 3.000 ;
        RECT  0.000 2.740 0.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.710 1.225 2.790 1.485 ;
        RECT  2.550 0.655 2.710 2.460 ;
        RECT  2.155 0.655 2.550 0.815 ;
        RECT  1.775 2.300 2.550 2.460 ;
        RECT  1.775 1.035 2.270 1.535 ;
        RECT  1.995 0.420 2.155 0.815 ;
        RECT  1.775 0.420 1.995 0.580 ;
        RECT  1.515 0.320 1.775 0.580 ;
        RECT  1.515 0.830 1.775 2.015 ;
        RECT  1.515 2.300 1.775 2.560 ;
        RECT  1.035 1.130 1.295 1.950 ;
        RECT  0.385 1.790 1.035 1.950 ;
        RECT  0.285 0.710 0.385 0.970 ;
        RECT  0.285 1.790 0.385 2.050 ;
        RECT  0.125 0.710 0.285 2.050 ;
    END
END DLY4X1MTH

MACRO DLY4X4MTH
    CLASS CORE ;
    FOREIGN DLY4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.930 1.045 4.000 1.730 ;
        RECT  3.670 0.610 3.930 1.730 ;
        RECT  3.455 1.570 3.670 1.730 ;
        RECT  3.195 1.570 3.455 2.435 ;
        END
        AntennaDiffArea 0.555 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 0.920 0.760 1.580 ;
        END
        AntennaGateArea 0.13 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 -0.130 4.100 0.130 ;
        RECT  3.100 -0.130 3.360 0.725 ;
        RECT  0.905 -0.130 3.100 0.130 ;
        RECT  0.645 -0.130 0.905 0.740 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 1.915 3.975 3.000 ;
        RECT  1.125 2.740 3.715 3.000 ;
        RECT  0.185 2.535 1.125 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.005 1.230 3.450 1.390 ;
        RECT  2.845 0.905 3.005 2.360 ;
        RECT  2.315 0.905 2.845 1.065 ;
        RECT  2.115 2.200 2.845 2.360 ;
        RECT  2.300 1.245 2.560 1.745 ;
        RECT  2.055 0.765 2.315 1.065 ;
        RECT  1.755 1.245 2.300 1.495 ;
        RECT  1.855 2.200 2.115 2.460 ;
        RECT  1.755 0.455 1.805 0.715 ;
        RECT  1.505 0.455 1.755 1.945 ;
        RECT  1.455 1.685 1.505 1.945 ;
        RECT  1.190 1.025 1.290 1.525 ;
        RECT  1.030 1.025 1.190 1.925 ;
        RECT  0.385 1.765 1.030 1.925 ;
        RECT  0.285 0.480 0.385 0.740 ;
        RECT  0.285 1.765 0.385 2.085 ;
        RECT  0.125 0.480 0.285 2.085 ;
    END
END DLY4X4MTH

MACRO EDFFHQX1MTH
    CLASS CORE ;
    FOREIGN EDFFHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.120 0.635 11.380 2.285 ;
        RECT  11.095 0.635 11.120 0.895 ;
        RECT  11.095 1.685 11.120 2.285 ;
        END
        AntennaDiffArea 0.34 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 0.705 1.635 1.540 ;
        RECT  1.290 1.225 1.475 1.540 ;
        END
        AntennaGateArea 0.1222 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.150 0.370 1.675 ;
        END
        AntennaGateArea 0.1209 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.415 0.920 4.450 1.170 ;
        RECT  4.020 0.680 4.415 1.170 ;
        RECT  3.950 1.010 4.020 1.170 ;
        END
        AntennaGateArea 0.1417 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.285 -0.130 11.480 0.130 ;
        RECT  11.025 -0.130 11.285 0.300 ;
        RECT  10.845 -0.130 11.025 0.130 ;
        RECT  10.585 -0.130 10.845 0.840 ;
        RECT  9.875 -0.130 10.585 0.300 ;
        RECT  7.595 -0.130 9.875 0.130 ;
        RECT  7.435 -0.130 7.595 0.300 ;
        RECT  3.055 -0.130 7.435 0.130 ;
        RECT  2.795 -0.130 3.055 0.300 ;
        RECT  1.450 -0.130 2.795 0.130 ;
        RECT  1.190 -0.130 1.450 0.300 ;
        RECT  0.725 -0.130 1.190 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 2.740 11.480 3.000 ;
        RECT  10.100 2.570 10.700 3.000 ;
        RECT  2.755 2.740 10.100 3.000 ;
        RECT  2.545 2.230 2.755 3.000 ;
        RECT  0.395 2.740 2.545 3.000 ;
        RECT  0.135 2.620 0.395 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.640 1.175 10.935 1.435 ;
        RECT  10.480 1.175 10.640 2.220 ;
        RECT  10.435 1.175 10.480 1.435 ;
        RECT  9.855 2.060 10.480 2.220 ;
        RECT  10.200 1.615 10.300 1.875 ;
        RECT  10.200 0.660 10.225 0.920 ;
        RECT  10.040 0.660 10.200 1.875 ;
        RECT  9.515 1.080 10.040 1.240 ;
        RECT  9.695 1.420 9.855 2.220 ;
        RECT  9.175 1.420 9.695 1.580 ;
        RECT  9.355 0.310 9.515 1.240 ;
        RECT  9.355 1.760 9.515 2.220 ;
        RECT  7.935 0.310 9.355 0.470 ;
        RECT  8.735 2.060 9.355 2.220 ;
        RECT  6.375 2.400 9.180 2.560 ;
        RECT  9.015 0.650 9.175 1.875 ;
        RECT  8.625 0.650 9.015 0.810 ;
        RECT  8.915 1.715 9.015 1.875 ;
        RECT  8.735 1.035 8.835 1.195 ;
        RECT  8.575 1.035 8.735 2.220 ;
        RECT  6.715 2.060 8.575 2.220 ;
        RECT  8.235 0.650 8.395 1.880 ;
        RECT  8.115 0.650 8.235 0.980 ;
        RECT  8.135 1.720 8.235 1.880 ;
        RECT  7.575 0.820 8.115 0.980 ;
        RECT  7.955 1.195 8.055 1.455 ;
        RECT  7.795 1.195 7.955 1.780 ;
        RECT  7.775 0.310 7.935 0.640 ;
        RECT  7.235 1.620 7.795 1.780 ;
        RECT  7.255 0.480 7.775 0.640 ;
        RECT  7.415 0.820 7.575 1.305 ;
        RECT  7.095 0.310 7.255 0.640 ;
        RECT  7.075 0.820 7.235 1.780 ;
        RECT  3.400 0.310 7.095 0.470 ;
        RECT  6.915 0.820 7.075 0.980 ;
        RECT  7.055 1.620 7.075 1.780 ;
        RECT  6.895 1.620 7.055 1.880 ;
        RECT  6.655 0.650 6.915 0.980 ;
        RECT  6.715 1.160 6.895 1.420 ;
        RECT  6.555 1.160 6.715 2.220 ;
        RECT  6.470 1.160 6.555 1.420 ;
        RECT  6.310 0.650 6.470 1.420 ;
        RECT  6.215 2.060 6.375 2.560 ;
        RECT  5.505 0.650 6.310 0.810 ;
        RECT  6.030 2.060 6.215 2.220 ;
        RECT  6.030 1.040 6.130 1.200 ;
        RECT  3.095 2.400 6.035 2.560 ;
        RECT  5.870 1.040 6.030 2.220 ;
        RECT  3.690 2.060 5.870 2.220 ;
        RECT  5.345 0.650 5.505 1.880 ;
        RECT  5.105 0.650 5.345 0.810 ;
        RECT  4.215 1.720 5.345 1.880 ;
        RECT  4.855 1.100 5.075 1.360 ;
        RECT  4.695 0.650 4.855 1.510 ;
        RECT  4.595 0.650 4.695 0.810 ;
        RECT  3.775 1.350 4.695 1.510 ;
        RECT  3.955 1.690 4.215 1.880 ;
        RECT  3.740 0.665 3.840 0.825 ;
        RECT  3.615 1.350 3.775 1.795 ;
        RECT  3.580 0.665 3.740 1.070 ;
        RECT  3.530 1.975 3.690 2.220 ;
        RECT  3.435 0.910 3.580 1.070 ;
        RECT  3.435 1.975 3.530 2.135 ;
        RECT  3.275 0.910 3.435 2.135 ;
        RECT  3.240 0.310 3.400 0.720 ;
        RECT  3.095 0.560 3.240 0.720 ;
        RECT  2.935 0.560 3.095 1.440 ;
        RECT  2.935 1.825 3.095 2.560 ;
        RECT  2.485 1.825 2.935 1.985 ;
        RECT  2.365 0.485 2.485 1.985 ;
        RECT  2.325 0.485 2.365 2.560 ;
        RECT  2.205 1.565 2.325 2.560 ;
        RECT  1.335 2.400 2.205 2.560 ;
        RECT  2.025 0.700 2.115 0.960 ;
        RECT  1.895 0.355 2.025 1.880 ;
        RECT  1.865 0.355 1.895 2.220 ;
        RECT  1.765 0.355 1.865 0.515 ;
        RECT  1.635 1.720 1.865 2.220 ;
        RECT  1.265 1.720 1.635 1.880 ;
        RECT  1.175 2.060 1.335 2.560 ;
        RECT  1.085 0.755 1.265 1.025 ;
        RECT  1.085 2.060 1.175 2.320 ;
        RECT  0.925 0.755 1.085 2.320 ;
        RECT  0.585 0.765 0.745 2.190 ;
    END
END EDFFHQX1MTH

MACRO EDFFHQX2MTH
    CLASS CORE ;
    FOREIGN EDFFHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.120 0.390 11.380 2.425 ;
        RECT  11.095 0.390 11.120 0.990 ;
        RECT  11.095 1.825 11.120 2.425 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 0.705 1.635 1.540 ;
        RECT  1.290 1.225 1.475 1.540 ;
        END
        AntennaGateArea 0.1248 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.150 0.370 1.675 ;
        END
        AntennaGateArea 0.0923 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.415 0.920 4.450 1.170 ;
        RECT  4.020 0.680 4.415 1.170 ;
        RECT  3.950 1.010 4.020 1.170 ;
        END
        AntennaGateArea 0.1443 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 -0.130 11.480 0.130 ;
        RECT  10.585 -0.130 10.845 0.840 ;
        RECT  9.875 -0.130 10.585 0.300 ;
        RECT  7.595 -0.130 9.875 0.130 ;
        RECT  7.435 -0.130 7.595 0.300 ;
        RECT  3.055 -0.130 7.435 0.130 ;
        RECT  2.795 -0.130 3.055 0.300 ;
        RECT  1.450 -0.130 2.795 0.130 ;
        RECT  1.190 -0.130 1.450 0.300 ;
        RECT  0.725 -0.130 1.190 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.700 2.740 11.480 3.000 ;
        RECT  10.100 2.570 10.700 3.000 ;
        RECT  2.755 2.740 10.100 3.000 ;
        RECT  2.545 2.230 2.755 3.000 ;
        RECT  0.385 2.740 2.545 3.000 ;
        RECT  0.125 2.620 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.575 1.205 10.935 1.465 ;
        RECT  10.415 1.205 10.575 2.220 ;
        RECT  9.855 2.060 10.415 2.220 ;
        RECT  10.205 0.660 10.265 0.920 ;
        RECT  10.045 0.660 10.205 1.875 ;
        RECT  9.515 1.080 10.045 1.240 ;
        RECT  9.695 1.420 9.855 2.220 ;
        RECT  9.175 1.420 9.695 1.580 ;
        RECT  9.355 0.310 9.515 1.240 ;
        RECT  9.355 1.760 9.515 2.220 ;
        RECT  7.935 0.310 9.355 0.470 ;
        RECT  8.735 2.060 9.355 2.220 ;
        RECT  6.375 2.400 9.180 2.560 ;
        RECT  9.015 0.650 9.175 1.875 ;
        RECT  8.625 0.650 9.015 0.810 ;
        RECT  8.915 1.715 9.015 1.875 ;
        RECT  8.735 1.035 8.835 1.195 ;
        RECT  8.575 1.035 8.735 2.220 ;
        RECT  6.715 2.060 8.575 2.220 ;
        RECT  8.235 0.650 8.395 1.880 ;
        RECT  8.115 0.650 8.235 0.980 ;
        RECT  8.135 1.720 8.235 1.880 ;
        RECT  7.575 0.820 8.115 0.980 ;
        RECT  7.955 1.195 8.055 1.455 ;
        RECT  7.795 1.195 7.955 1.780 ;
        RECT  7.775 0.310 7.935 0.640 ;
        RECT  7.235 1.620 7.795 1.780 ;
        RECT  7.255 0.480 7.775 0.640 ;
        RECT  7.415 0.820 7.575 1.305 ;
        RECT  7.095 0.310 7.255 0.640 ;
        RECT  7.075 0.820 7.235 1.780 ;
        RECT  3.400 0.310 7.095 0.470 ;
        RECT  6.915 0.820 7.075 0.980 ;
        RECT  7.055 1.620 7.075 1.780 ;
        RECT  6.895 1.620 7.055 1.880 ;
        RECT  6.655 0.650 6.915 0.980 ;
        RECT  6.715 1.160 6.895 1.420 ;
        RECT  6.555 1.160 6.715 2.220 ;
        RECT  6.470 1.160 6.555 1.420 ;
        RECT  6.310 0.650 6.470 1.420 ;
        RECT  6.215 2.060 6.375 2.560 ;
        RECT  5.505 0.650 6.310 0.810 ;
        RECT  6.030 2.060 6.215 2.220 ;
        RECT  6.030 0.990 6.130 1.150 ;
        RECT  3.095 2.400 6.035 2.560 ;
        RECT  5.870 0.990 6.030 2.220 ;
        RECT  3.690 2.060 5.870 2.220 ;
        RECT  5.345 0.650 5.505 1.875 ;
        RECT  5.105 0.650 5.345 0.810 ;
        RECT  4.355 1.715 5.345 1.875 ;
        RECT  4.855 1.100 5.075 1.360 ;
        RECT  4.695 0.650 4.855 1.510 ;
        RECT  4.595 0.650 4.695 0.810 ;
        RECT  3.845 1.350 4.695 1.510 ;
        RECT  4.095 1.690 4.355 1.875 ;
        RECT  3.685 1.350 3.845 1.795 ;
        RECT  3.740 0.665 3.840 0.825 ;
        RECT  3.580 0.665 3.740 1.070 ;
        RECT  3.530 1.975 3.690 2.220 ;
        RECT  3.615 1.535 3.685 1.795 ;
        RECT  3.435 0.910 3.580 1.070 ;
        RECT  3.435 1.975 3.530 2.135 ;
        RECT  3.275 0.910 3.435 2.135 ;
        RECT  3.240 0.310 3.400 0.720 ;
        RECT  3.095 0.560 3.240 0.720 ;
        RECT  2.935 0.560 3.095 1.440 ;
        RECT  2.935 1.825 3.095 2.560 ;
        RECT  2.485 1.825 2.935 1.985 ;
        RECT  2.365 0.485 2.485 1.985 ;
        RECT  2.325 0.485 2.365 2.560 ;
        RECT  2.205 1.565 2.325 2.560 ;
        RECT  1.335 2.400 2.205 2.560 ;
        RECT  2.025 0.700 2.115 0.960 ;
        RECT  1.895 0.355 2.025 1.880 ;
        RECT  1.865 0.355 1.895 2.220 ;
        RECT  1.765 0.355 1.865 0.515 ;
        RECT  1.635 1.720 1.865 2.220 ;
        RECT  1.275 1.720 1.635 1.880 ;
        RECT  1.175 2.130 1.335 2.560 ;
        RECT  1.095 0.755 1.265 1.015 ;
        RECT  1.095 2.130 1.175 2.390 ;
        RECT  0.935 0.755 1.095 2.390 ;
        RECT  0.585 0.755 0.745 2.190 ;
    END
END EDFFHQX2MTH

MACRO EDFFHQX4MTH
    CLASS CORE ;
    FOREIGN EDFFHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.665 1.290 11.790 1.580 ;
        RECT  11.405 0.390 11.665 2.425 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.685 2.045 1.355 ;
        END
        AntennaGateArea 0.13 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.275 1.285 0.720 1.705 ;
        END
        AntennaGateArea 0.1651 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.825 0.920 4.860 1.170 ;
        RECT  4.445 0.680 4.825 1.170 ;
        RECT  4.360 1.010 4.445 1.170 ;
        END
        AntennaGateArea 0.1859 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 -0.130 12.300 0.130 ;
        RECT  11.915 -0.130 12.175 0.990 ;
        RECT  11.125 -0.130 11.915 0.130 ;
        RECT  10.525 -0.130 11.125 0.300 ;
        RECT  8.055 -0.130 10.525 0.130 ;
        RECT  7.895 -0.130 8.055 0.300 ;
        RECT  3.465 -0.130 7.895 0.130 ;
        RECT  3.205 -0.130 3.465 0.300 ;
        RECT  1.865 -0.130 3.205 0.130 ;
        RECT  1.265 -0.130 1.865 0.300 ;
        RECT  0.560 -0.130 1.265 0.130 ;
        RECT  0.300 -0.130 0.560 0.980 ;
        RECT  0.000 -0.130 0.300 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 2.740 12.300 3.000 ;
        RECT  11.915 1.825 12.175 3.000 ;
        RECT  11.125 2.740 11.915 3.000 ;
        RECT  10.525 2.570 11.125 3.000 ;
        RECT  3.645 2.740 10.525 3.000 ;
        RECT  3.045 2.620 3.645 3.000 ;
        RECT  0.525 2.740 3.045 3.000 ;
        RECT  0.265 1.890 0.525 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.915 1.205 11.075 2.365 ;
        RECT  10.305 2.205 10.915 2.365 ;
        RECT  10.485 0.765 10.645 1.945 ;
        RECT  10.275 0.765 10.485 0.925 ;
        RECT  10.145 1.420 10.305 2.365 ;
        RECT  10.115 0.310 10.275 1.195 ;
        RECT  9.895 1.420 10.145 1.580 ;
        RECT  8.395 0.310 10.115 0.470 ;
        RECT  9.795 1.760 9.955 2.220 ;
        RECT  9.735 0.650 9.895 1.580 ;
        RECT  9.145 2.060 9.795 2.220 ;
        RECT  9.015 0.650 9.735 0.810 ;
        RECT  9.585 1.420 9.735 1.580 ;
        RECT  9.425 1.420 9.585 1.875 ;
        RECT  6.785 2.400 9.575 2.560 ;
        RECT  9.145 1.020 9.535 1.180 ;
        RECT  9.325 1.715 9.425 1.875 ;
        RECT  8.985 1.020 9.145 2.220 ;
        RECT  7.125 2.060 8.985 2.220 ;
        RECT  8.645 0.745 8.805 1.880 ;
        RECT  8.555 0.745 8.645 1.005 ;
        RECT  8.545 1.720 8.645 1.880 ;
        RECT  7.985 0.845 8.555 1.005 ;
        RECT  8.365 1.195 8.465 1.455 ;
        RECT  8.235 0.310 8.395 0.640 ;
        RECT  8.205 1.195 8.365 1.780 ;
        RECT  7.665 0.480 8.235 0.640 ;
        RECT  7.645 1.620 8.205 1.780 ;
        RECT  7.825 0.845 7.985 1.375 ;
        RECT  7.505 0.310 7.665 0.640 ;
        RECT  7.485 0.820 7.645 1.780 ;
        RECT  3.810 0.310 7.505 0.470 ;
        RECT  7.325 0.820 7.485 0.980 ;
        RECT  7.465 1.620 7.485 1.780 ;
        RECT  7.305 1.620 7.465 1.880 ;
        RECT  7.065 0.650 7.325 0.980 ;
        RECT  7.125 1.160 7.305 1.420 ;
        RECT  6.965 1.160 7.125 2.220 ;
        RECT  6.880 1.160 6.965 1.420 ;
        RECT  6.720 0.650 6.880 1.420 ;
        RECT  6.625 2.060 6.785 2.560 ;
        RECT  5.915 0.650 6.720 0.810 ;
        RECT  6.440 2.060 6.625 2.220 ;
        RECT  6.440 0.990 6.540 1.150 ;
        RECT  3.985 2.400 6.445 2.560 ;
        RECT  6.280 0.990 6.440 2.220 ;
        RECT  4.325 2.060 6.280 2.220 ;
        RECT  5.755 0.650 5.915 1.875 ;
        RECT  5.515 0.650 5.755 0.810 ;
        RECT  4.765 1.715 5.755 1.875 ;
        RECT  5.265 1.180 5.485 1.440 ;
        RECT  5.105 0.650 5.265 1.510 ;
        RECT  5.005 0.650 5.105 0.810 ;
        RECT  4.235 1.350 5.105 1.510 ;
        RECT  4.505 1.690 4.765 1.875 ;
        RECT  4.165 1.925 4.325 2.220 ;
        RECT  4.165 0.650 4.265 0.810 ;
        RECT  4.075 1.350 4.235 1.730 ;
        RECT  4.005 0.650 4.165 1.070 ;
        RECT  3.795 1.925 4.165 2.085 ;
        RECT  3.975 1.570 4.075 1.730 ;
        RECT  3.795 0.910 4.005 1.070 ;
        RECT  3.825 2.270 3.985 2.560 ;
        RECT  2.735 2.270 3.825 2.430 ;
        RECT  3.650 0.310 3.810 0.720 ;
        RECT  3.635 0.910 3.795 2.085 ;
        RECT  3.455 0.560 3.650 0.720 ;
        RECT  3.295 0.560 3.455 1.460 ;
        RECT  3.255 1.200 3.295 1.460 ;
        RECT  2.835 0.520 2.995 1.730 ;
        RECT  2.735 0.520 2.835 0.780 ;
        RECT  2.735 1.570 2.835 1.730 ;
        RECT  2.575 1.570 2.735 2.560 ;
        RECT  1.575 2.400 2.575 2.560 ;
        RECT  2.385 0.720 2.525 0.980 ;
        RECT  2.225 0.310 2.385 1.720 ;
        RECT  2.115 1.560 2.225 1.720 ;
        RECT  2.115 2.060 2.215 2.220 ;
        RECT  1.955 1.560 2.115 2.220 ;
        RECT  1.705 1.560 1.955 1.720 ;
        RECT  1.525 1.890 1.575 2.560 ;
        RECT  1.525 0.745 1.560 1.005 ;
        RECT  1.365 0.745 1.525 2.560 ;
        RECT  1.315 1.890 1.365 2.560 ;
        RECT  1.065 0.745 1.100 1.005 ;
        RECT  0.905 0.745 1.065 2.490 ;
        RECT  0.840 0.745 0.905 1.005 ;
        RECT  0.805 1.890 0.905 2.490 ;
    END
END EDFFHQX4MTH

MACRO EDFFHQX8MTH
    CLASS CORE ;
    FOREIGN EDFFHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.635 0.390 12.895 2.425 ;
        RECT  11.875 1.170 12.635 1.735 ;
        RECT  11.615 0.390 11.875 2.425 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.170 2.360 1.785 ;
        END
        AntennaGateArea 0.1313 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.275 1.285 0.720 1.705 ;
        END
        AntennaGateArea 0.1651 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.740 0.880 4.820 1.170 ;
        RECT  4.435 0.680 4.740 1.170 ;
        RECT  4.350 1.010 4.435 1.170 ;
        END
        AntennaGateArea 0.1859 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 -0.130 13.530 0.130 ;
        RECT  13.145 -0.130 13.405 0.990 ;
        RECT  12.385 -0.130 13.145 0.130 ;
        RECT  12.125 -0.130 12.385 0.990 ;
        RECT  11.365 -0.130 12.125 0.130 ;
        RECT  11.105 -0.130 11.365 0.990 ;
        RECT  10.525 -0.130 11.105 0.300 ;
        RECT  8.045 -0.130 10.525 0.130 ;
        RECT  7.885 -0.130 8.045 0.300 ;
        RECT  3.460 -0.130 7.885 0.130 ;
        RECT  3.200 -0.130 3.460 0.300 ;
        RECT  1.495 -0.130 3.200 0.130 ;
        RECT  1.235 -0.130 1.495 0.300 ;
        RECT  0.400 -0.130 1.235 0.130 ;
        RECT  0.140 -0.130 0.400 0.980 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.825 13.405 3.000 ;
        RECT  12.385 2.740 13.145 3.000 ;
        RECT  12.125 1.915 12.385 3.000 ;
        RECT  11.395 2.740 12.125 3.000 ;
        RECT  11.155 1.760 11.395 3.000 ;
        RECT  10.430 2.565 11.155 3.000 ;
        RECT  3.625 2.740 10.430 3.000 ;
        RECT  3.025 2.620 3.625 3.000 ;
        RECT  0.510 2.740 3.025 3.000 ;
        RECT  0.250 1.890 0.510 3.000 ;
        RECT  0.000 2.740 0.250 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.975 1.205 11.355 1.465 ;
        RECT  10.815 1.205 10.975 2.285 ;
        RECT  10.285 2.125 10.815 2.285 ;
        RECT  10.635 0.765 10.735 1.025 ;
        RECT  10.485 0.765 10.635 1.945 ;
        RECT  10.475 0.595 10.485 1.945 ;
        RECT  10.265 0.595 10.475 1.195 ;
        RECT  10.125 1.420 10.285 2.285 ;
        RECT  10.105 0.310 10.265 1.195 ;
        RECT  9.885 1.420 10.125 1.580 ;
        RECT  8.385 0.310 10.105 0.470 ;
        RECT  9.785 1.760 9.945 2.220 ;
        RECT  9.725 0.650 9.885 1.580 ;
        RECT  9.135 2.060 9.785 2.220 ;
        RECT  9.005 0.650 9.725 0.810 ;
        RECT  9.575 1.420 9.725 1.580 ;
        RECT  9.415 1.420 9.575 1.875 ;
        RECT  6.775 2.400 9.565 2.560 ;
        RECT  9.135 1.020 9.525 1.180 ;
        RECT  9.315 1.715 9.415 1.875 ;
        RECT  8.975 1.020 9.135 2.220 ;
        RECT  7.115 2.060 8.975 2.220 ;
        RECT  8.635 0.745 8.795 1.880 ;
        RECT  8.545 0.745 8.635 1.005 ;
        RECT  8.535 1.720 8.635 1.880 ;
        RECT  7.975 0.820 8.545 0.980 ;
        RECT  8.355 1.195 8.455 1.455 ;
        RECT  8.225 0.310 8.385 0.640 ;
        RECT  8.195 1.195 8.355 1.780 ;
        RECT  7.655 0.480 8.225 0.640 ;
        RECT  7.635 1.620 8.195 1.780 ;
        RECT  7.815 0.820 7.975 1.375 ;
        RECT  7.495 0.310 7.655 0.640 ;
        RECT  7.475 0.820 7.635 1.780 ;
        RECT  3.800 0.310 7.495 0.470 ;
        RECT  7.315 0.820 7.475 0.980 ;
        RECT  7.455 1.620 7.475 1.780 ;
        RECT  7.295 1.620 7.455 1.880 ;
        RECT  7.055 0.650 7.315 0.980 ;
        RECT  7.115 1.160 7.295 1.420 ;
        RECT  6.955 1.160 7.115 2.220 ;
        RECT  6.870 1.160 6.955 1.420 ;
        RECT  6.710 0.650 6.870 1.420 ;
        RECT  6.615 2.060 6.775 2.560 ;
        RECT  5.905 0.650 6.710 0.810 ;
        RECT  6.430 2.060 6.615 2.220 ;
        RECT  6.430 0.990 6.530 1.150 ;
        RECT  3.975 2.400 6.435 2.560 ;
        RECT  6.270 0.990 6.430 2.220 ;
        RECT  4.315 2.060 6.270 2.220 ;
        RECT  5.745 0.650 5.905 1.875 ;
        RECT  5.505 0.650 5.745 0.810 ;
        RECT  4.755 1.715 5.745 1.875 ;
        RECT  5.255 1.180 5.475 1.440 ;
        RECT  5.095 0.650 5.255 1.510 ;
        RECT  4.995 0.650 5.095 0.810 ;
        RECT  4.225 1.350 5.095 1.510 ;
        RECT  4.495 1.690 4.755 1.875 ;
        RECT  4.155 1.925 4.315 2.220 ;
        RECT  4.155 0.650 4.255 0.810 ;
        RECT  4.065 1.350 4.225 1.730 ;
        RECT  3.995 0.650 4.155 1.070 ;
        RECT  3.785 1.925 4.155 2.085 ;
        RECT  3.965 1.570 4.065 1.730 ;
        RECT  3.785 0.910 3.995 1.070 ;
        RECT  3.815 2.270 3.975 2.560 ;
        RECT  2.700 2.270 3.815 2.430 ;
        RECT  3.640 0.310 3.800 0.720 ;
        RECT  3.625 0.910 3.785 2.085 ;
        RECT  3.395 0.560 3.640 0.720 ;
        RECT  3.235 0.560 3.395 1.265 ;
        RECT  2.015 0.310 2.965 0.470 ;
        RECT  2.540 0.650 2.700 2.560 ;
        RECT  2.345 0.650 2.540 0.810 ;
        RECT  1.560 2.400 2.540 2.560 ;
        RECT  1.905 2.060 2.165 2.220 ;
        RECT  1.905 0.310 2.015 0.615 ;
        RECT  1.745 0.310 1.905 2.220 ;
        RECT  1.590 1.485 1.745 1.745 ;
        RECT  1.400 1.940 1.560 2.560 ;
        RECT  1.240 0.745 1.400 2.560 ;
        RECT  0.900 0.745 1.060 2.490 ;
        RECT  0.680 0.745 0.900 1.005 ;
        RECT  0.790 1.890 0.900 2.490 ;
    END
END EDFFHQX8MTH

MACRO EDFFTRX1MTH
    CLASS CORE ;
    FOREIGN EDFFTRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.220 1.270 4.860 1.540 ;
        END
        AntennaGateArea 0.052 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.160 1.700 12.200 1.990 ;
        RECT  12.155 1.700 12.160 2.320 ;
        RECT  11.995 0.715 12.155 2.320 ;
        RECT  11.965 0.715 11.995 0.975 ;
        RECT  11.900 1.700 11.995 2.320 ;
        END
        AntennaDiffArea 0.34 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.090 0.835 11.380 1.170 ;
        RECT  10.930 0.835 11.090 2.320 ;
        RECT  10.900 0.835 10.930 0.995 ;
        END
        AntennaDiffArea 0.349 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 0.920 3.630 1.130 ;
        RECT  3.305 0.920 3.465 1.540 ;
        RECT  1.400 1.380 3.305 1.540 ;
        RECT  1.240 1.200 1.400 1.540 ;
        END
        AntennaGateArea 0.1066 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.810 1.125 4.040 1.540 ;
        RECT  3.645 1.330 3.810 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.375 1.720 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.965 -0.130 12.300 0.130 ;
        RECT  11.025 -0.130 11.965 0.290 ;
        RECT  6.500 -0.130 11.025 0.130 ;
        RECT  6.240 -0.130 6.500 0.760 ;
        RECT  4.715 -0.130 6.240 0.130 ;
        RECT  4.555 -0.130 4.715 0.485 ;
        RECT  1.155 -0.130 4.555 0.130 ;
        RECT  0.555 -0.130 1.155 0.470 ;
        RECT  0.000 -0.130 0.555 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.650 2.740 12.300 3.000 ;
        RECT  11.390 1.720 11.650 3.000 ;
        RECT  10.450 2.740 11.390 3.000 ;
        RECT  9.950 2.300 10.450 3.000 ;
        RECT  1.525 2.740 9.950 3.000 ;
        RECT  0.585 2.500 1.525 3.000 ;
        RECT  0.000 2.740 0.585 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.785 1.235 11.815 1.495 ;
        RECT  11.625 0.475 11.785 1.495 ;
        RECT  10.750 0.475 11.625 0.635 ;
        RECT  10.720 0.355 10.750 0.635 ;
        RECT  10.560 0.355 10.720 1.960 ;
        RECT  10.490 0.355 10.560 0.515 ;
        RECT  9.770 1.800 10.560 1.960 ;
        RECT  10.310 1.050 10.380 1.310 ;
        RECT  10.150 0.395 10.310 1.310 ;
        RECT  9.090 0.395 10.150 0.555 ;
        RECT  9.610 1.390 9.770 2.560 ;
        RECT  9.430 0.880 9.630 1.040 ;
        RECT  2.170 2.400 9.610 2.560 ;
        RECT  9.270 0.880 9.430 2.220 ;
        RECT  7.910 2.060 9.270 2.220 ;
        RECT  8.930 0.395 9.090 1.880 ;
        RECT  8.770 0.395 8.930 0.555 ;
        RECT  8.690 1.720 8.930 1.880 ;
        RECT  8.510 0.870 8.750 1.030 ;
        RECT  7.910 1.350 8.750 1.510 ;
        RECT  8.350 0.375 8.510 1.030 ;
        RECT  7.540 0.375 8.350 0.535 ;
        RECT  7.750 0.715 7.910 2.220 ;
        RECT  5.220 2.060 7.750 2.220 ;
        RECT  7.540 1.720 7.570 1.880 ;
        RECT  7.380 0.375 7.540 1.880 ;
        RECT  6.920 0.375 7.380 0.535 ;
        RECT  7.310 1.720 7.380 1.880 ;
        RECT  7.070 1.195 7.200 1.455 ;
        RECT  6.910 0.790 7.070 1.880 ;
        RECT  6.810 0.790 6.910 1.100 ;
        RECT  6.800 1.720 6.910 1.880 ;
        RECT  6.290 0.940 6.810 1.100 ;
        RECT  6.560 1.280 6.720 1.540 ;
        RECT  6.220 1.380 6.560 1.540 ;
        RECT  6.030 0.940 6.290 1.200 ;
        RECT  6.060 1.380 6.220 1.850 ;
        RECT  5.560 1.690 6.060 1.850 ;
        RECT  5.400 0.620 5.560 1.850 ;
        RECT  5.060 0.430 5.220 2.220 ;
        RECT  4.925 0.430 5.060 0.690 ;
        RECT  1.645 1.720 5.060 1.880 ;
        RECT  4.555 0.785 4.715 1.060 ;
        RECT  1.985 2.060 4.685 2.220 ;
        RECT  4.095 0.785 4.555 0.945 ;
        RECT  3.935 0.475 4.095 0.945 ;
        RECT  2.085 0.475 3.935 0.635 ;
        RECT  2.775 0.815 3.035 1.055 ;
        RECT  1.055 0.815 2.775 0.975 ;
        RECT  1.825 2.060 1.985 2.320 ;
        RECT  1.485 1.720 1.645 2.320 ;
        RECT  0.715 2.160 1.485 2.320 ;
        RECT  1.145 1.720 1.305 1.980 ;
        RECT  1.055 1.720 1.145 1.880 ;
        RECT  0.895 0.815 1.055 1.880 ;
        RECT  0.555 0.865 0.715 2.320 ;
        RECT  0.340 0.865 0.555 1.025 ;
        RECT  0.125 1.900 0.555 2.060 ;
        RECT  0.180 0.765 0.340 1.025 ;
    END
END EDFFTRX1MTH

MACRO EDFFTRX2MTH
    CLASS CORE ;
    FOREIGN EDFFTRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.390 1.270 4.860 1.540 ;
        END
        AntennaGateArea 0.052 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.525 1.290 12.610 1.580 ;
        RECT  12.365 0.425 12.525 2.320 ;
        RECT  12.245 1.720 12.365 2.320 ;
        END
        AntennaDiffArea 0.548 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.480 1.250 11.790 1.580 ;
        RECT  11.480 0.815 11.585 0.975 ;
        RECT  11.220 0.815 11.480 2.320 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.880 3.590 1.540 ;
        RECT  1.400 1.380 3.380 1.540 ;
        RECT  1.240 1.200 1.400 1.540 ;
        END
        AntennaGateArea 0.1066 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.165 4.050 1.425 ;
        RECT  3.785 0.880 4.000 1.425 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.375 1.720 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.505 -0.130 12.710 0.130 ;
        RECT  9.905 -0.130 10.505 0.250 ;
        RECT  6.625 -0.130 9.905 0.130 ;
        RECT  6.365 -0.130 6.625 0.870 ;
        RECT  5.300 -0.130 6.365 0.130 ;
        RECT  4.700 -0.130 5.300 0.325 ;
        RECT  1.640 -0.130 4.700 0.130 ;
        RECT  0.700 -0.130 1.640 0.515 ;
        RECT  0.000 -0.130 0.700 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.995 2.740 12.710 3.000 ;
        RECT  11.735 1.890 11.995 3.000 ;
        RECT  10.790 2.740 11.735 3.000 ;
        RECT  10.290 2.370 10.790 3.000 ;
        RECT  1.610 2.740 10.290 3.000 ;
        RECT  0.670 2.435 1.610 3.000 ;
        RECT  0.000 2.740 0.670 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.025 0.475 12.185 1.495 ;
        RECT  11.025 0.475 12.025 0.635 ;
        RECT  10.865 0.450 11.025 1.960 ;
        RECT  10.110 1.800 10.865 1.960 ;
        RECT  10.525 0.440 10.685 1.440 ;
        RECT  9.655 0.440 10.525 0.600 ;
        RECT  9.950 1.345 10.110 2.560 ;
        RECT  2.270 2.400 9.950 2.560 ;
        RECT  9.765 0.880 9.935 1.040 ;
        RECT  9.605 0.880 9.765 2.220 ;
        RECT  9.425 0.410 9.655 0.600 ;
        RECT  8.230 2.060 9.605 2.220 ;
        RECT  9.265 0.410 9.425 1.880 ;
        RECT  9.055 0.410 9.265 0.600 ;
        RECT  9.100 1.720 9.265 1.880 ;
        RECT  8.825 0.870 9.085 1.030 ;
        RECT  8.230 1.350 9.085 1.510 ;
        RECT  8.665 0.415 8.825 1.030 ;
        RECT  7.720 0.415 8.665 0.575 ;
        RECT  8.070 0.765 8.230 2.220 ;
        RECT  7.915 0.765 8.070 0.925 ;
        RECT  5.300 2.060 8.070 2.220 ;
        RECT  7.720 1.720 7.890 1.880 ;
        RECT  7.560 0.415 7.720 1.880 ;
        RECT  7.100 0.415 7.560 0.575 ;
        RECT  7.290 1.195 7.380 1.455 ;
        RECT  7.290 1.720 7.320 1.880 ;
        RECT  7.130 0.800 7.290 1.880 ;
        RECT  6.990 0.800 7.130 1.210 ;
        RECT  7.060 1.720 7.130 1.880 ;
        RECT  6.460 1.050 6.990 1.210 ;
        RECT  6.825 1.390 6.950 1.550 ;
        RECT  6.665 1.390 6.825 1.845 ;
        RECT  5.645 1.685 6.665 1.845 ;
        RECT  6.200 1.050 6.460 1.260 ;
        RECT  5.485 0.730 5.645 1.845 ;
        RECT  5.385 0.730 5.485 0.890 ;
        RECT  5.140 1.170 5.300 2.220 ;
        RECT  5.060 1.170 5.140 1.880 ;
        RECT  1.750 1.720 5.060 1.880 ;
        RECT  4.340 0.850 4.970 1.010 ;
        RECT  2.090 2.060 4.960 2.220 ;
        RECT  4.180 0.520 4.340 1.010 ;
        RECT  2.165 0.520 4.180 0.680 ;
        RECT  1.740 0.895 3.130 1.055 ;
        RECT  1.930 2.060 2.090 2.320 ;
        RECT  1.590 1.720 1.750 2.235 ;
        RECT  1.580 0.815 1.740 1.055 ;
        RECT  0.715 2.075 1.590 2.235 ;
        RECT  1.055 0.815 1.580 0.975 ;
        RECT  1.055 1.735 1.410 1.895 ;
        RECT  0.895 0.815 1.055 1.895 ;
        RECT  0.555 0.865 0.715 2.235 ;
        RECT  0.340 0.865 0.555 1.025 ;
        RECT  0.125 1.900 0.555 2.060 ;
        RECT  0.180 0.765 0.340 1.025 ;
    END
END EDFFTRX2MTH

MACRO EDFFTRX4MTH
    CLASS CORE ;
    FOREIGN EDFFTRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.940 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.330 1.270 4.860 1.540 ;
        END
        AntennaGateArea 0.052 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.315 1.290 13.430 1.580 ;
        RECT  13.155 0.425 13.315 2.320 ;
        RECT  13.095 0.425 13.155 1.025 ;
        RECT  13.045 1.720 13.155 2.320 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.115 0.815 12.375 2.320 ;
        RECT  11.990 1.250 12.115 1.580 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.880 3.590 1.540 ;
        RECT  1.840 1.380 3.380 1.540 ;
        RECT  1.240 1.280 1.840 1.540 ;
        END
        AntennaGateArea 0.1066 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.165 4.050 1.425 ;
        RECT  3.785 0.880 4.000 1.425 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.375 1.720 ;
        END
        AntennaGateArea 0.1053 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.815 -0.130 13.940 0.130 ;
        RECT  13.555 -0.130 13.815 0.985 ;
        RECT  11.835 -0.130 13.555 0.130 ;
        RECT  11.575 -0.130 11.835 0.290 ;
        RECT  10.810 -0.130 11.575 0.130 ;
        RECT  10.210 -0.130 10.810 0.250 ;
        RECT  8.340 -0.130 10.210 0.130 ;
        RECT  8.080 -0.130 8.340 0.250 ;
        RECT  6.560 -0.130 8.080 0.130 ;
        RECT  6.300 -0.130 6.560 0.810 ;
        RECT  5.300 -0.130 6.300 0.130 ;
        RECT  4.700 -0.130 5.300 0.350 ;
        RECT  1.640 -0.130 4.700 0.130 ;
        RECT  0.700 -0.130 1.640 0.515 ;
        RECT  0.000 -0.130 0.700 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.760 2.740 13.940 3.000 ;
        RECT  13.760 1.815 13.815 2.415 ;
        RECT  13.600 1.815 13.760 3.000 ;
        RECT  13.555 1.815 13.600 2.415 ;
        RECT  11.815 2.740 13.600 3.000 ;
        RECT  11.655 1.895 11.815 3.000 ;
        RECT  10.760 2.740 11.655 3.000 ;
        RECT  10.600 2.485 10.760 3.000 ;
        RECT  1.610 2.740 10.600 3.000 ;
        RECT  0.670 2.520 1.610 3.000 ;
        RECT  0.000 2.740 0.670 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.910 1.235 12.975 1.495 ;
        RECT  12.750 0.475 12.910 1.495 ;
        RECT  11.475 0.475 12.750 0.635 ;
        RECT  11.350 0.475 11.475 2.180 ;
        RECT  11.315 0.475 11.350 2.380 ;
        RECT  11.090 0.475 11.315 0.785 ;
        RECT  11.090 1.880 11.315 2.380 ;
        RECT  10.970 0.970 11.130 1.700 ;
        RECT  10.420 2.020 11.090 2.180 ;
        RECT  10.525 0.970 10.970 1.130 ;
        RECT  10.365 0.490 10.525 1.130 ;
        RECT  10.260 1.450 10.420 2.560 ;
        RECT  9.740 0.490 10.365 0.650 ;
        RECT  2.270 2.400 10.260 2.560 ;
        RECT  9.920 0.970 10.080 2.220 ;
        RECT  8.235 2.060 9.920 2.220 ;
        RECT  9.580 0.490 9.740 1.880 ;
        RECT  9.175 0.490 9.580 0.650 ;
        RECT  9.210 1.720 9.580 1.880 ;
        RECT  9.240 0.885 9.400 1.145 ;
        RECT  8.965 0.985 9.240 1.145 ;
        RECT  8.235 1.415 9.085 1.575 ;
        RECT  8.805 0.430 8.965 1.145 ;
        RECT  7.720 0.430 8.805 0.590 ;
        RECT  8.075 0.770 8.235 2.220 ;
        RECT  7.900 0.770 8.075 1.030 ;
        RECT  5.300 2.060 8.075 2.220 ;
        RECT  7.720 1.690 7.850 1.850 ;
        RECT  7.560 0.310 7.720 1.850 ;
        RECT  7.015 0.310 7.560 0.470 ;
        RECT  7.340 1.250 7.380 1.510 ;
        RECT  7.290 1.250 7.340 1.850 ;
        RECT  7.150 0.970 7.290 1.850 ;
        RECT  7.130 0.680 7.150 1.850 ;
        RECT  6.890 0.680 7.130 1.155 ;
        RECT  7.080 1.690 7.130 1.850 ;
        RECT  6.825 1.335 6.950 1.495 ;
        RECT  6.465 0.995 6.890 1.155 ;
        RECT  6.665 1.335 6.825 1.845 ;
        RECT  5.645 1.685 6.665 1.845 ;
        RECT  6.205 0.995 6.465 1.210 ;
        RECT  5.485 0.730 5.645 1.845 ;
        RECT  5.385 0.730 5.485 0.890 ;
        RECT  5.140 1.130 5.300 2.220 ;
        RECT  5.060 1.130 5.140 1.880 ;
        RECT  1.750 1.720 5.060 1.880 ;
        RECT  4.345 0.790 4.960 0.950 ;
        RECT  2.090 2.060 4.960 2.220 ;
        RECT  4.340 0.520 4.345 0.950 ;
        RECT  4.180 0.520 4.340 1.000 ;
        RECT  2.165 0.520 4.180 0.680 ;
        RECT  1.985 0.895 3.130 1.055 ;
        RECT  1.930 2.060 2.090 2.320 ;
        RECT  1.825 0.815 1.985 1.055 ;
        RECT  1.055 0.815 1.825 0.975 ;
        RECT  1.590 1.720 1.750 2.235 ;
        RECT  0.715 2.075 1.590 2.235 ;
        RECT  1.055 1.735 1.410 1.895 ;
        RECT  0.895 0.815 1.055 1.895 ;
        RECT  0.555 0.865 0.715 2.235 ;
        RECT  0.340 0.865 0.555 1.025 ;
        RECT  0.125 1.900 0.555 2.060 ;
        RECT  0.180 0.765 0.340 1.025 ;
    END
END EDFFTRX4MTH

MACRO EDFFX1MTH
    CLASS CORE ;
    FOREIGN EDFFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.050 0.735 11.310 1.990 ;
        RECT  10.760 1.700 11.050 1.990 ;
        END
        AntennaDiffArea 0.348 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.205 0.735 10.270 0.995 ;
        RECT  9.945 0.735 10.205 1.955 ;
        RECT  9.940 1.290 9.945 1.580 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.200 1.855 1.360 ;
        RECT  0.445 1.200 0.720 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.220 2.815 1.480 ;
        RECT  2.560 0.880 2.770 1.480 ;
        RECT  2.555 1.220 2.560 1.480 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.300 1.280 5.790 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.125 -0.130 11.480 0.130 ;
        RECT  10.780 -0.130 11.125 0.300 ;
        RECT  10.520 -0.130 10.780 0.995 ;
        RECT  10.185 -0.130 10.520 0.300 ;
        RECT  9.840 -0.130 10.185 0.130 ;
        RECT  8.900 -0.130 9.840 0.300 ;
        RECT  5.830 -0.130 8.900 0.130 ;
        RECT  5.670 -0.130 5.830 0.300 ;
        RECT  0.745 -0.130 5.670 0.130 ;
        RECT  0.145 -0.130 0.745 0.300 ;
        RECT  0.000 -0.130 0.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.745 2.740 11.480 3.000 ;
        RECT  10.485 2.475 10.745 3.000 ;
        RECT  9.985 2.740 10.485 3.000 ;
        RECT  9.045 2.570 9.985 3.000 ;
        RECT  3.825 2.740 9.045 3.000 ;
        RECT  3.225 2.620 3.825 3.000 ;
        RECT  2.780 2.740 3.225 3.000 ;
        RECT  1.840 2.620 2.780 3.000 ;
        RECT  1.065 2.740 1.840 3.000 ;
        RECT  0.725 2.570 1.065 3.000 ;
        RECT  0.125 2.285 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.710 1.200 10.870 1.460 ;
        RECT  10.560 1.300 10.710 1.460 ;
        RECT  10.400 1.300 10.560 2.295 ;
        RECT  9.730 2.135 10.400 2.295 ;
        RECT  9.730 0.765 9.760 1.025 ;
        RECT  9.570 0.765 9.730 2.295 ;
        RECT  9.500 0.765 9.570 1.025 ;
        RECT  9.380 1.810 9.570 2.070 ;
        RECT  9.230 1.245 9.390 1.505 ;
        RECT  8.815 1.860 9.380 2.020 ;
        RECT  8.390 1.250 9.230 1.410 ;
        RECT  8.655 1.860 8.815 2.560 ;
        RECT  4.245 2.400 8.655 2.560 ;
        RECT  8.045 0.310 8.640 0.470 ;
        RECT  8.385 0.715 8.390 1.410 ;
        RECT  8.250 0.715 8.385 2.045 ;
        RECT  8.230 0.715 8.250 2.220 ;
        RECT  8.225 1.250 8.230 2.220 ;
        RECT  8.090 1.885 8.225 2.220 ;
        RECT  7.910 0.310 8.045 1.705 ;
        RECT  7.885 0.310 7.910 2.220 ;
        RECT  6.170 0.310 7.885 0.470 ;
        RECT  7.750 1.545 7.885 2.220 ;
        RECT  4.590 2.060 7.750 2.220 ;
        RECT  7.570 1.085 7.705 1.345 ;
        RECT  7.410 0.940 7.570 1.850 ;
        RECT  6.645 0.940 7.410 1.100 ;
        RECT  6.310 1.690 7.410 1.850 ;
        RECT  6.130 1.320 7.230 1.480 ;
        RECT  6.385 0.650 6.645 1.100 ;
        RECT  5.485 0.940 6.385 1.100 ;
        RECT  6.010 0.310 6.170 0.760 ;
        RECT  5.970 1.320 6.130 1.880 ;
        RECT  5.875 0.480 6.010 0.760 ;
        RECT  5.120 1.720 5.970 1.880 ;
        RECT  5.325 0.310 5.485 1.100 ;
        RECT  3.985 0.310 5.325 0.470 ;
        RECT  5.120 0.650 5.145 0.910 ;
        RECT  4.960 0.650 5.120 1.880 ;
        RECT  4.465 0.650 4.960 0.810 ;
        RECT  4.770 1.720 4.960 1.880 ;
        RECT  4.620 1.205 4.780 1.540 ;
        RECT  3.645 1.380 4.620 1.540 ;
        RECT  4.430 1.940 4.590 2.220 ;
        RECT  4.305 0.650 4.465 0.985 ;
        RECT  3.275 1.940 4.430 2.100 ;
        RECT  4.085 2.280 4.245 2.560 ;
        RECT  1.535 2.280 4.085 2.440 ;
        RECT  3.825 0.310 3.985 1.170 ;
        RECT  3.485 0.455 3.645 1.760 ;
        RECT  3.115 0.790 3.275 2.100 ;
        RECT  1.065 0.380 3.125 0.540 ;
        RECT  3.015 0.790 3.115 0.950 ;
        RECT  2.775 1.840 2.935 2.100 ;
        RECT  1.065 1.895 2.775 2.055 ;
        RECT  2.235 1.510 2.335 1.670 ;
        RECT  2.075 0.720 2.235 1.670 ;
        RECT  1.685 0.720 2.075 0.880 ;
        RECT  1.525 0.720 1.685 0.975 ;
        RECT  1.275 2.280 1.535 2.505 ;
        RECT  0.265 0.815 1.525 0.975 ;
        RECT  0.555 1.760 0.815 2.020 ;
        RECT  0.265 1.760 0.555 1.920 ;
        RECT  0.105 0.815 0.265 1.920 ;
    END
END EDFFX1MTH

MACRO EDFFX2MTH
    CLASS CORE ;
    FOREIGN EDFFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.050 0.425 11.310 2.285 ;
        RECT  10.760 1.700 11.050 1.990 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.205 0.425 10.270 1.025 ;
        RECT  9.940 0.425 10.205 1.945 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.200 1.850 1.360 ;
        RECT  0.445 1.200 0.720 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.220 2.815 1.480 ;
        RECT  2.555 0.880 2.770 1.480 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 1.280 5.765 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.780 -0.130 11.480 0.130 ;
        RECT  10.520 -0.130 10.780 0.975 ;
        RECT  9.660 -0.130 10.520 0.130 ;
        RECT  8.820 -0.130 9.660 0.300 ;
        RECT  7.670 -0.130 8.820 0.130 ;
        RECT  7.170 -0.130 7.670 0.300 ;
        RECT  5.830 -0.130 7.170 0.130 ;
        RECT  5.670 -0.130 5.830 0.300 ;
        RECT  0.815 -0.130 5.670 0.130 ;
        RECT  0.215 -0.130 0.815 0.505 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.745 2.740 11.480 3.000 ;
        RECT  10.485 2.570 10.745 3.000 ;
        RECT  9.670 2.740 10.485 3.000 ;
        RECT  9.070 2.570 9.670 3.000 ;
        RECT  3.690 2.740 9.070 3.000 ;
        RECT  3.090 2.620 3.690 3.000 ;
        RECT  2.735 2.740 3.090 3.000 ;
        RECT  1.795 2.620 2.735 3.000 ;
        RECT  1.065 2.740 1.795 3.000 ;
        RECT  0.725 2.570 1.065 3.000 ;
        RECT  0.125 2.285 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.710 1.200 10.870 1.460 ;
        RECT  10.560 1.300 10.710 1.460 ;
        RECT  10.400 1.300 10.560 2.295 ;
        RECT  9.730 2.135 10.400 2.295 ;
        RECT  9.730 0.765 9.760 1.025 ;
        RECT  9.570 0.765 9.730 2.295 ;
        RECT  9.500 0.765 9.570 1.025 ;
        RECT  9.430 1.810 9.570 2.070 ;
        RECT  8.890 1.860 9.430 2.020 ;
        RECT  9.230 1.245 9.390 1.505 ;
        RECT  8.480 1.245 9.230 1.405 ;
        RECT  8.730 1.860 8.890 2.560 ;
        RECT  4.180 2.400 8.730 2.560 ;
        RECT  8.050 0.310 8.640 0.470 ;
        RECT  8.390 1.245 8.480 2.185 ;
        RECT  8.320 0.715 8.390 2.185 ;
        RECT  8.230 0.715 8.320 1.405 ;
        RECT  8.090 2.025 8.320 2.185 ;
        RECT  8.050 1.645 8.140 1.805 ;
        RECT  7.910 0.310 8.050 1.805 ;
        RECT  7.890 0.310 7.910 2.220 ;
        RECT  6.990 0.600 7.890 0.760 ;
        RECT  7.750 1.645 7.890 2.220 ;
        RECT  4.525 2.060 7.750 2.220 ;
        RECT  7.570 1.115 7.710 1.375 ;
        RECT  7.410 0.940 7.570 1.850 ;
        RECT  6.650 0.940 7.410 1.100 ;
        RECT  6.315 1.690 7.410 1.850 ;
        RECT  6.105 1.320 7.230 1.480 ;
        RECT  6.830 0.310 6.990 0.760 ;
        RECT  6.210 0.310 6.830 0.470 ;
        RECT  6.390 0.650 6.650 1.100 ;
        RECT  5.485 0.940 6.390 1.100 ;
        RECT  6.050 0.310 6.210 0.760 ;
        RECT  5.945 1.320 6.105 1.880 ;
        RECT  5.875 0.600 6.050 0.760 ;
        RECT  5.115 1.720 5.945 1.880 ;
        RECT  5.325 0.310 5.485 1.100 ;
        RECT  3.985 0.310 5.325 0.470 ;
        RECT  5.115 0.650 5.145 0.940 ;
        RECT  4.955 0.650 5.115 1.880 ;
        RECT  4.465 0.650 4.955 0.810 ;
        RECT  4.770 1.650 4.955 1.880 ;
        RECT  4.615 1.205 4.775 1.465 ;
        RECT  4.325 1.305 4.615 1.465 ;
        RECT  4.365 1.940 4.525 2.220 ;
        RECT  4.305 0.650 4.465 0.985 ;
        RECT  3.305 1.940 4.365 2.100 ;
        RECT  4.165 1.305 4.325 1.540 ;
        RECT  4.020 2.280 4.180 2.560 ;
        RECT  3.645 1.380 4.165 1.540 ;
        RECT  1.505 2.280 4.020 2.440 ;
        RECT  3.825 0.310 3.985 1.130 ;
        RECT  3.485 0.450 3.645 1.760 ;
        RECT  3.145 0.790 3.305 2.100 ;
        RECT  3.015 0.790 3.145 0.950 ;
        RECT  1.065 0.380 3.125 0.540 ;
        RECT  2.805 1.745 2.965 2.055 ;
        RECT  1.065 1.895 2.805 2.055 ;
        RECT  2.235 1.510 2.335 1.670 ;
        RECT  2.075 0.720 2.235 1.670 ;
        RECT  1.685 0.720 2.075 0.880 ;
        RECT  1.525 0.720 1.685 0.975 ;
        RECT  0.265 0.815 1.525 0.975 ;
        RECT  1.245 2.280 1.505 2.550 ;
        RECT  0.555 1.760 0.815 2.020 ;
        RECT  0.265 1.760 0.555 1.920 ;
        RECT  0.105 0.815 0.265 1.920 ;
    END
END EDFFX2MTH

MACRO EDFFX4MTH
    CLASS CORE ;
    FOREIGN EDFFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.420 0.425 11.680 2.295 ;
        RECT  11.400 1.695 11.420 2.295 ;
        RECT  11.170 1.695 11.400 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.570 0.425 10.640 1.025 ;
        RECT  10.310 0.425 10.570 1.955 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.200 1.855 1.360 ;
        RECT  0.445 1.200 0.720 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.220 2.815 1.480 ;
        RECT  2.555 0.880 2.770 1.480 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.295 1.280 5.790 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.170 -0.130 12.300 0.130 ;
        RECT  11.910 -0.130 12.170 0.955 ;
        RECT  11.150 -0.130 11.910 0.130 ;
        RECT  10.890 -0.130 11.150 0.975 ;
        RECT  10.010 -0.130 10.890 0.130 ;
        RECT  9.070 -0.130 10.010 0.300 ;
        RECT  5.845 -0.130 9.070 0.130 ;
        RECT  5.685 -0.130 5.845 0.300 ;
        RECT  0.725 -0.130 5.685 0.130 ;
        RECT  0.125 -0.130 0.725 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.170 2.740 12.300 3.000 ;
        RECT  11.910 1.915 12.170 3.000 ;
        RECT  11.115 2.740 11.910 3.000 ;
        RECT  10.855 2.570 11.115 3.000 ;
        RECT  10.020 2.740 10.855 3.000 ;
        RECT  9.080 2.570 10.020 3.000 ;
        RECT  3.890 2.740 9.080 3.000 ;
        RECT  2.950 2.620 3.890 3.000 ;
        RECT  2.645 2.740 2.950 3.000 ;
        RECT  1.705 2.620 2.645 3.000 ;
        RECT  1.065 2.740 1.705 3.000 ;
        RECT  0.725 2.570 1.065 3.000 ;
        RECT  0.125 2.285 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.080 1.200 11.240 1.460 ;
        RECT  10.910 1.300 11.080 1.460 ;
        RECT  10.750 1.300 10.910 2.295 ;
        RECT  10.130 2.135 10.750 2.295 ;
        RECT  9.970 0.865 10.130 2.295 ;
        RECT  9.730 0.865 9.970 1.025 ;
        RECT  9.400 1.900 9.970 2.160 ;
        RECT  9.280 1.245 9.790 1.505 ;
        RECT  9.470 0.765 9.730 1.025 ;
        RECT  8.885 2.000 9.400 2.160 ;
        RECT  8.480 1.245 9.280 1.405 ;
        RECT  8.725 2.000 8.885 2.560 ;
        RECT  4.250 2.400 8.725 2.560 ;
        RECT  8.045 0.310 8.640 0.470 ;
        RECT  8.320 0.715 8.480 2.185 ;
        RECT  8.230 0.715 8.320 0.975 ;
        RECT  8.100 2.025 8.320 2.185 ;
        RECT  8.045 1.645 8.140 1.805 ;
        RECT  7.910 0.310 8.045 1.805 ;
        RECT  7.885 0.310 7.910 2.220 ;
        RECT  6.205 0.310 7.885 0.470 ;
        RECT  7.750 1.645 7.885 2.220 ;
        RECT  4.590 2.060 7.750 2.220 ;
        RECT  7.570 1.105 7.705 1.365 ;
        RECT  7.410 0.940 7.570 1.850 ;
        RECT  6.645 0.940 7.410 1.100 ;
        RECT  6.310 1.690 7.410 1.850 ;
        RECT  6.130 1.320 7.230 1.480 ;
        RECT  6.385 0.650 6.645 1.100 ;
        RECT  5.505 0.940 6.385 1.100 ;
        RECT  6.045 0.310 6.205 0.760 ;
        RECT  5.970 1.320 6.130 1.880 ;
        RECT  5.875 0.540 6.045 0.760 ;
        RECT  5.115 1.720 5.970 1.880 ;
        RECT  5.345 0.310 5.505 1.100 ;
        RECT  3.985 0.310 5.345 0.470 ;
        RECT  5.115 0.650 5.165 0.910 ;
        RECT  4.955 0.650 5.115 1.880 ;
        RECT  4.465 0.650 4.955 0.810 ;
        RECT  4.770 1.720 4.955 1.880 ;
        RECT  4.615 1.205 4.775 1.540 ;
        RECT  3.645 1.380 4.615 1.540 ;
        RECT  4.430 1.940 4.590 2.220 ;
        RECT  4.305 0.650 4.465 0.985 ;
        RECT  3.305 1.940 4.430 2.100 ;
        RECT  4.090 2.280 4.250 2.560 ;
        RECT  1.505 2.280 4.090 2.440 ;
        RECT  3.825 0.310 3.985 1.170 ;
        RECT  3.485 0.455 3.645 1.760 ;
        RECT  3.145 0.790 3.305 2.100 ;
        RECT  3.015 0.790 3.145 0.950 ;
        RECT  1.065 0.380 3.125 0.540 ;
        RECT  2.805 1.745 2.965 2.055 ;
        RECT  1.065 1.895 2.805 2.055 ;
        RECT  2.235 1.510 2.335 1.670 ;
        RECT  2.075 0.720 2.235 1.670 ;
        RECT  1.685 0.720 2.075 0.880 ;
        RECT  1.525 0.720 1.685 0.975 ;
        RECT  0.265 0.815 1.525 0.975 ;
        RECT  1.245 2.280 1.505 2.500 ;
        RECT  0.555 1.760 0.815 2.020 ;
        RECT  0.265 1.760 0.555 1.920 ;
        RECT  0.105 0.815 0.265 1.920 ;
    END
END EDFFX4MTH

MACRO FILL16MTH
    CLASS CORE SPACER ;
    FOREIGN FILL16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 6.560 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 6.560 3.000 ;
        END
    END VDD
END FILL16MTH

MACRO FILL1MTH
    CLASS CORE SPACER ;
    FOREIGN FILL1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.410 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 0.410 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 0.410 3.000 ;
        END
    END VDD
END FILL1MTH

MACRO FILL2MTH
    CLASS CORE SPACER ;
    FOREIGN FILL2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.820 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 0.820 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 0.820 3.000 ;
        END
    END VDD
END FILL2MTH

MACRO FILL32MTH
    CLASS CORE SPACER ;
    FOREIGN FILL32MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.120 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 13.120 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 13.120 3.000 ;
        END
    END VDD
END FILL32MTH

MACRO FILL4MTH
    CLASS CORE SPACER ;
    FOREIGN FILL4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 1.640 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 1.640 3.000 ;
        END
    END VDD
END FILL4MTH

MACRO FILL64MTH
    CLASS CORE SPACER ;
    FOREIGN FILL64MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.240 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 26.240 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 26.240 3.000 ;
        END
    END VDD
END FILL64MTH

MACRO FILL8MTH
    CLASS CORE SPACER ;
    FOREIGN FILL8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 -0.130 3.280 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.000 2.740 3.280 3.000 ;
        END
    END VDD
END FILL8MTH

MACRO FILLCAP16MTH
    CLASS CORE SPACER ;
    FOREIGN FILLCAP16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.980 ;
        RECT  0.000 -0.130 6.175 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 6.560 3.000 ;
        RECT  0.125 1.850 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.275 1.185 6.415 1.345 ;
        RECT  6.115 1.185 6.275 2.410 ;
        RECT  6.015 1.785 6.115 2.410 ;
        RECT  0.335 0.405 0.495 1.525 ;
        RECT  0.145 1.365 0.335 1.525 ;
    END
END FILLCAP16MTH

MACRO FILLCAP32MTH
    CLASS CORE SPACER ;
    FOREIGN FILLCAP32MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.120 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.995 -0.130 13.120 0.130 ;
        RECT  12.735 -0.130 12.995 0.980 ;
        RECT  0.000 -0.130 12.735 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 13.120 3.000 ;
        RECT  0.125 1.850 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.835 1.185 12.975 1.345 ;
        RECT  12.675 1.185 12.835 2.410 ;
        RECT  12.575 1.785 12.675 2.410 ;
        RECT  0.335 0.405 0.495 1.525 ;
        RECT  0.145 1.365 0.335 1.525 ;
    END
END FILLCAP32MTH

MACRO FILLCAP4MTH
    CLASS CORE SPACER ;
    FOREIGN FILLCAP4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.515 -0.130 1.640 0.130 ;
        RECT  1.255 -0.130 1.515 0.980 ;
        RECT  0.000 -0.130 1.255 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 1.640 3.000 ;
        RECT  0.125 1.850 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.355 1.185 1.495 1.345 ;
        RECT  1.195 1.185 1.355 2.410 ;
        RECT  1.095 1.785 1.195 2.410 ;
        RECT  0.335 0.405 0.495 1.525 ;
        RECT  0.145 1.365 0.335 1.525 ;
    END
END FILLCAP4MTH

MACRO FILLCAP64MTH
    CLASS CORE SPACER ;
    FOREIGN FILLCAP64MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 26.240 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  26.115 -0.130 26.240 0.130 ;
        RECT  25.855 -0.130 26.115 0.980 ;
        RECT  0.000 -0.130 25.855 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 26.240 3.000 ;
        RECT  0.125 1.850 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  25.955 1.185 26.095 1.345 ;
        RECT  25.795 1.185 25.955 2.410 ;
        RECT  25.695 1.785 25.795 2.410 ;
        RECT  0.335 0.405 0.495 1.525 ;
        RECT  0.145 1.365 0.335 1.525 ;
    END
END FILLCAP64MTH

MACRO FILLCAP8MTH
    CLASS CORE SPACER ;
    FOREIGN FILLCAP8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 -0.130 3.280 0.130 ;
        RECT  2.895 -0.130 3.155 0.980 ;
        RECT  0.000 -0.130 2.895 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 3.280 3.000 ;
        RECT  0.125 1.850 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.995 1.185 3.135 1.345 ;
        RECT  2.835 1.185 2.995 2.410 ;
        RECT  2.735 1.785 2.835 2.410 ;
        RECT  0.335 0.405 0.495 1.525 ;
        RECT  0.145 1.365 0.335 1.525 ;
    END
END FILLCAP8MTH

MACRO FILLTIEMTH
    CLASS CORE ;
    FOREIGN FILLTIEMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.820 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 -0.130 0.820 0.130 ;
        RECT  0.280 -0.130 0.540 0.995 ;
        RECT  0.000 -0.130 0.280 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 2.740 0.820 3.000 ;
        RECT  0.280 1.805 0.540 3.000 ;
        RECT  0.000 2.740 0.280 3.000 ;
        END
    END VDD
END FILLTIEMTH

MACRO HOLDX1MTH
    CLASS CORE ;
    FOREIGN HOLDX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION INOUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.355 0.365 1.515 1.990 ;
        RECT  1.245 0.365 1.355 0.625 ;
        RECT  0.920 1.580 1.355 1.990 ;
        RECT  0.745 1.580 0.920 1.740 ;
        RECT  0.585 1.135 0.745 1.740 ;
        RECT  0.440 1.135 0.585 1.395 ;
        END
        AntennaGateArea 0.0533 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 -0.130 1.640 0.130 ;
        RECT  0.645 -0.130 0.905 0.300 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.965 2.740 1.640 3.000 ;
        RECT  0.705 2.230 0.965 3.000 ;
        RECT  0.000 2.740 0.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.925 0.795 1.085 1.400 ;
        RECT  0.385 0.795 0.925 0.955 ;
        RECT  0.260 0.335 0.385 0.955 ;
        RECT  0.260 1.685 0.385 1.945 ;
        RECT  0.100 0.335 0.260 1.945 ;
    END
END HOLDX1MTH

MACRO INVX10MTH
    CLASS CORE ;
    FOREIGN INVX10MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 0.410 3.085 2.420 ;
        RECT  2.065 1.085 2.825 1.785 ;
        RECT  1.805 0.405 2.065 2.420 ;
        RECT  1.430 0.795 1.805 2.075 ;
        RECT  1.045 0.795 1.430 1.110 ;
        RECT  1.045 1.720 1.430 2.075 ;
        RECT  0.785 0.410 1.045 1.110 ;
        RECT  0.785 1.720 1.045 2.420 ;
        END
        AntennaDiffArea 1.737 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.290 1.215 1.540 ;
        END
        AntennaGateArea 1.027 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 -0.130 3.280 0.130 ;
        RECT  2.315 -0.130 2.575 0.905 ;
        RECT  1.555 -0.130 2.315 0.130 ;
        RECT  1.295 -0.130 1.555 0.615 ;
        RECT  0.505 -0.130 1.295 0.130 ;
        RECT  0.245 -0.130 0.505 0.980 ;
        RECT  0.000 -0.130 0.245 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 2.740 3.280 3.000 ;
        RECT  2.315 1.965 2.575 3.000 ;
        RECT  1.555 2.740 2.315 3.000 ;
        RECT  1.295 2.255 1.555 3.000 ;
        RECT  0.505 2.740 1.295 3.000 ;
        RECT  0.245 1.890 0.505 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
END INVX10MTH

MACRO INVX12MTH
    CLASS CORE ;
    FOREIGN INVX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.715 0.410 2.975 2.385 ;
        RECT  1.955 1.085 2.715 1.785 ;
        RECT  1.695 0.405 1.955 2.420 ;
        RECT  0.935 0.745 1.695 1.095 ;
        RECT  0.935 1.725 1.695 2.125 ;
        RECT  0.675 0.410 0.935 1.095 ;
        RECT  0.675 1.725 0.935 2.420 ;
        END
        AntennaDiffArea 1.8 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.280 1.445 1.540 ;
        END
        AntennaGateArea 1.2324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 -0.130 3.690 0.130 ;
        RECT  3.265 -0.130 3.525 1.010 ;
        RECT  2.465 -0.130 3.265 0.130 ;
        RECT  2.205 -0.130 2.465 0.905 ;
        RECT  1.445 -0.130 2.205 0.130 ;
        RECT  1.185 -0.130 1.445 0.565 ;
        RECT  0.385 -0.130 1.185 0.130 ;
        RECT  0.125 -0.130 0.385 1.010 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 2.740 3.690 3.000 ;
        RECT  3.265 1.780 3.525 3.000 ;
        RECT  2.465 2.740 3.265 3.000 ;
        RECT  2.205 1.965 2.465 3.000 ;
        RECT  1.445 2.740 2.205 3.000 ;
        RECT  1.185 2.305 1.445 3.000 ;
        RECT  0.385 2.740 1.185 3.000 ;
        RECT  0.125 1.780 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX12MTH

MACRO INVX14MTH
    CLASS CORE ;
    FOREIGN INVX14MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 0.410 3.955 2.420 ;
        RECT  2.935 0.745 3.695 1.745 ;
        RECT  2.675 0.410 2.935 2.420 ;
        RECT  1.915 0.745 2.675 1.745 ;
        RECT  1.655 0.405 1.915 2.420 ;
        RECT  1.260 0.745 1.655 2.125 ;
        RECT  0.925 0.745 1.260 1.125 ;
        RECT  0.925 1.745 1.260 2.125 ;
        RECT  0.605 0.410 0.925 1.125 ;
        RECT  0.605 1.745 0.925 2.420 ;
        END
        AntennaDiffArea 2.337 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.305 1.075 1.565 ;
        END
        AntennaGateArea 1.4378 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 -0.130 4.100 0.130 ;
        RECT  3.185 -0.130 3.445 0.565 ;
        RECT  2.425 -0.130 3.185 0.130 ;
        RECT  2.165 -0.130 2.425 0.565 ;
        RECT  1.405 -0.130 2.165 0.130 ;
        RECT  1.145 -0.130 1.405 0.565 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.985 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 2.740 4.100 3.000 ;
        RECT  3.185 1.965 3.445 3.000 ;
        RECT  2.425 2.740 3.185 3.000 ;
        RECT  2.165 1.960 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 2.305 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.915 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX14MTH

MACRO INVX16MTH
    CLASS CORE ;
    FOREIGN INVX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 0.410 3.875 2.420 ;
        RECT  2.935 1.085 3.615 1.785 ;
        RECT  2.675 0.410 2.935 2.420 ;
        RECT  1.915 1.085 2.675 1.785 ;
        RECT  1.655 0.405 1.915 2.420 ;
        RECT  1.585 0.745 1.655 2.125 ;
        RECT  0.895 0.745 1.585 1.140 ;
        RECT  0.895 1.720 1.585 2.125 ;
        RECT  0.635 0.410 0.895 1.140 ;
        RECT  0.635 1.720 0.895 2.420 ;
        END
        AntennaDiffArea 2.4 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.320 1.405 1.540 ;
        END
        AntennaGateArea 1.6432 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  4.125 -0.130 4.385 0.955 ;
        RECT  2.425 -0.130 4.125 0.130 ;
        RECT  2.165 -0.130 2.425 0.905 ;
        RECT  1.405 -0.130 2.165 0.130 ;
        RECT  1.145 -0.130 1.405 0.565 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 1.010 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.915 4.385 3.000 ;
        RECT  2.425 2.740 4.125 3.000 ;
        RECT  2.165 1.965 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 2.305 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.780 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX16MTH

MACRO INVX18MTH
    CLASS CORE ;
    FOREIGN INVX18MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.535 0.410 4.795 1.075 ;
        RECT  4.535 1.755 4.795 2.355 ;
        RECT  3.775 0.745 4.535 1.075 ;
        RECT  3.775 1.755 4.535 2.075 ;
        RECT  3.515 0.410 3.775 2.360 ;
        RECT  2.785 0.745 3.515 2.075 ;
        RECT  2.350 0.420 2.785 2.385 ;
        RECT  0.635 0.420 2.350 1.075 ;
        RECT  0.635 1.785 2.350 2.385 ;
        END
        AntennaDiffArea 2.937 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 1.300 1.745 1.540 ;
        END
        AntennaGateArea 1.8486 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 -0.130 4.920 0.130 ;
        RECT  4.025 -0.130 4.285 0.565 ;
        RECT  3.265 -0.130 4.025 0.130 ;
        RECT  3.005 -0.130 3.265 0.565 ;
        RECT  0.385 -0.130 3.005 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 2.740 4.920 3.000 ;
        RECT  4.025 2.255 4.285 3.000 ;
        RECT  3.265 2.740 4.025 3.000 ;
        RECT  3.005 2.255 3.265 3.000 ;
        RECT  0.385 2.740 3.005 3.000 ;
        RECT  0.125 1.860 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX18MTH

MACRO INVX1MTH
    CLASS CORE ;
    FOREIGN INVX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.750 1.130 2.020 ;
        RECT  0.650 0.750 0.920 1.010 ;
        RECT  0.650 1.760 0.920 2.020 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.190 0.720 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 -0.130 1.230 0.130 ;
        RECT  0.400 -0.130 1.080 0.300 ;
        RECT  0.140 -0.130 0.400 0.970 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.080 2.740 1.230 3.000 ;
        RECT  0.400 2.570 1.080 3.000 ;
        RECT  0.140 1.825 0.400 3.000 ;
        RECT  0.000 2.740 0.140 3.000 ;
        END
    END VDD
END INVX1MTH

MACRO INVX20MTH
    CLASS CORE ;
    FOREIGN INVX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.780 0.410 5.040 1.110 ;
        RECT  4.780 1.720 5.040 2.360 ;
        RECT  4.020 0.745 4.780 1.110 ;
        RECT  4.020 1.720 4.780 2.125 ;
        RECT  3.760 0.410 4.020 2.360 ;
        RECT  3.000 0.745 3.760 2.125 ;
        RECT  2.740 0.405 3.000 2.360 ;
        RECT  2.420 0.745 2.740 2.125 ;
        RECT  2.015 0.745 2.420 1.110 ;
        RECT  1.980 1.720 2.420 2.125 ;
        RECT  1.720 0.410 2.015 1.110 ;
        RECT  1.720 1.720 1.980 2.360 ;
        RECT  0.960 0.745 1.720 1.110 ;
        RECT  0.960 1.720 1.720 2.125 ;
        RECT  0.700 0.410 0.960 1.110 ;
        RECT  0.700 1.720 0.960 2.360 ;
        END
        AntennaDiffArea 3 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.530 1.290 1.470 1.540 ;
        RECT  0.470 1.330 0.530 1.540 ;
        END
        AntennaGateArea 2.054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.580 -0.130 5.740 0.130 ;
        RECT  5.320 -0.130 5.580 0.980 ;
        RECT  4.530 -0.130 5.320 0.130 ;
        RECT  4.270 -0.130 4.530 0.565 ;
        RECT  3.510 -0.130 4.270 0.130 ;
        RECT  3.250 -0.130 3.510 0.565 ;
        RECT  2.490 -0.130 3.250 0.130 ;
        RECT  2.230 -0.130 2.490 0.565 ;
        RECT  1.470 -0.130 2.230 0.130 ;
        RECT  1.210 -0.130 1.470 0.565 ;
        RECT  0.420 -0.130 1.210 0.130 ;
        RECT  0.160 -0.130 0.420 0.980 ;
        RECT  0.000 -0.130 0.160 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.580 2.740 5.740 3.000 ;
        RECT  5.320 1.890 5.580 3.000 ;
        RECT  4.530 2.740 5.320 3.000 ;
        RECT  4.270 2.305 4.530 3.000 ;
        RECT  3.510 2.740 4.270 3.000 ;
        RECT  3.250 2.305 3.510 3.000 ;
        RECT  2.490 2.740 3.250 3.000 ;
        RECT  2.230 2.305 2.490 3.000 ;
        RECT  1.470 2.740 2.230 3.000 ;
        RECT  1.210 2.305 1.470 3.000 ;
        RECT  0.420 2.740 1.210 3.000 ;
        RECT  0.160 1.890 0.420 3.000 ;
        RECT  0.000 2.740 0.160 3.000 ;
        END
    END VDD
END INVX20MTH

MACRO INVX24MTH
    CLASS CORE ;
    FOREIGN INVX24MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.665 0.410 5.925 2.420 ;
        RECT  4.975 1.085 5.665 1.785 ;
        RECT  4.715 0.405 4.975 2.420 ;
        RECT  3.955 1.085 4.715 1.785 ;
        RECT  3.695 0.410 3.955 2.420 ;
        RECT  2.935 1.085 3.695 1.785 ;
        RECT  2.675 0.410 2.935 2.420 ;
        RECT  1.915 1.085 2.675 1.785 ;
        RECT  1.655 0.405 1.915 2.420 ;
        RECT  0.895 0.835 1.655 1.095 ;
        RECT  0.895 1.720 1.655 1.980 ;
        RECT  0.635 0.410 0.895 1.095 ;
        RECT  0.635 1.720 0.895 2.420 ;
        END
        AntennaDiffArea 3.6 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.275 1.405 1.540 ;
        END
        AntennaGateArea 2.4648 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.955 ;
        RECT  4.465 -0.130 6.175 0.130 ;
        RECT  4.205 -0.130 4.465 0.905 ;
        RECT  3.445 -0.130 4.205 0.130 ;
        RECT  3.185 -0.130 3.445 0.905 ;
        RECT  2.425 -0.130 3.185 0.130 ;
        RECT  2.165 -0.130 2.425 0.905 ;
        RECT  1.405 -0.130 2.165 0.130 ;
        RECT  1.145 -0.130 1.405 0.655 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 1.010 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.915 6.435 3.000 ;
        RECT  4.465 2.740 6.175 3.000 ;
        RECT  4.205 1.965 4.465 3.000 ;
        RECT  3.445 2.740 4.205 3.000 ;
        RECT  3.185 1.965 3.445 3.000 ;
        RECT  2.425 2.740 3.185 3.000 ;
        RECT  2.165 1.965 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 2.160 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.780 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX24MTH

MACRO INVX2MTH
    CLASS CORE ;
    FOREIGN INVX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 0.795 1.130 1.990 ;
        RECT  0.920 0.795 0.950 2.410 ;
        RECT  0.650 0.405 0.920 1.005 ;
        RECT  0.690 1.760 0.920 2.410 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.190 0.720 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 -0.130 1.230 0.130 ;
        RECT  0.140 -0.130 0.400 0.980 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 2.740 1.230 3.000 ;
        RECT  0.140 1.850 0.400 3.000 ;
        RECT  0.000 2.740 0.140 3.000 ;
        END
    END VDD
END INVX2MTH

MACRO INVX32MTH
    CLASS CORE ;
    FOREIGN INVX32MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.715 0.410 7.975 2.420 ;
        RECT  7.015 1.125 7.715 1.745 ;
        RECT  6.755 0.410 7.015 2.420 ;
        RECT  5.995 1.125 6.755 1.745 ;
        RECT  5.735 0.405 5.995 2.420 ;
        RECT  4.975 1.125 5.735 1.745 ;
        RECT  4.715 0.410 4.975 2.420 ;
        RECT  3.955 1.125 4.715 1.745 ;
        RECT  3.695 0.410 3.955 2.420 ;
        RECT  2.935 1.125 3.695 1.745 ;
        RECT  2.675 0.410 2.935 2.420 ;
        RECT  1.915 1.125 2.675 1.745 ;
        RECT  1.655 0.405 1.915 2.420 ;
        RECT  0.895 0.840 1.655 1.100 ;
        RECT  0.895 1.720 1.655 1.980 ;
        RECT  0.635 0.410 0.895 1.100 ;
        RECT  0.635 1.720 0.895 2.420 ;
        END
        AntennaDiffArea 4.8 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.280 1.405 1.540 ;
        END
        AntennaGateArea 3.2864 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.485 -0.130 8.610 0.130 ;
        RECT  8.225 -0.130 8.485 0.955 ;
        RECT  6.505 -0.130 8.225 0.130 ;
        RECT  6.245 -0.130 6.505 0.905 ;
        RECT  5.485 -0.130 6.245 0.130 ;
        RECT  5.225 -0.130 5.485 0.905 ;
        RECT  4.465 -0.130 5.225 0.130 ;
        RECT  4.205 -0.130 4.465 0.905 ;
        RECT  3.445 -0.130 4.205 0.130 ;
        RECT  3.185 -0.130 3.445 0.905 ;
        RECT  2.425 -0.130 3.185 0.130 ;
        RECT  2.165 -0.130 2.425 0.905 ;
        RECT  1.405 -0.130 2.165 0.130 ;
        RECT  1.145 -0.130 1.405 0.660 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.485 2.740 8.610 3.000 ;
        RECT  8.225 1.925 8.485 3.000 ;
        RECT  6.505 2.740 8.225 3.000 ;
        RECT  6.245 1.925 6.505 3.000 ;
        RECT  5.485 2.740 6.245 3.000 ;
        RECT  5.225 1.925 5.485 3.000 ;
        RECT  4.465 2.740 5.225 3.000 ;
        RECT  4.205 1.925 4.465 3.000 ;
        RECT  3.445 2.740 4.205 3.000 ;
        RECT  3.185 1.925 3.445 3.000 ;
        RECT  2.425 2.740 3.185 3.000 ;
        RECT  2.165 1.925 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 2.160 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.915 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX32MTH

MACRO INVX3MTH
    CLASS CORE ;
    FOREIGN INVX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.880 1.540 1.990 ;
        RECT  0.935 0.880 1.330 1.040 ;
        RECT  0.935 1.765 1.330 1.990 ;
        RECT  0.680 0.580 0.935 1.040 ;
        RECT  0.675 1.765 0.935 2.365 ;
        END
        AntennaDiffArea 0.456 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.505 1.290 1.105 1.580 ;
        END
        AntennaGateArea 0.312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 -0.130 1.640 0.130 ;
        RECT  1.225 -0.130 1.485 0.700 ;
        RECT  0.385 -0.130 1.225 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 2.740 1.640 3.000 ;
        RECT  1.225 2.170 1.485 3.000 ;
        RECT  0.385 2.740 1.225 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX3MTH

MACRO INVX4MTH
    CLASS CORE ;
    FOREIGN INVX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.880 1.540 1.990 ;
        RECT  0.935 0.880 1.330 1.040 ;
        RECT  0.935 1.765 1.330 1.990 ;
        RECT  0.680 0.580 0.935 1.040 ;
        RECT  0.680 1.765 0.935 2.365 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.505 1.290 1.105 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 -0.130 1.640 0.130 ;
        RECT  1.225 -0.130 1.485 0.700 ;
        RECT  0.385 -0.130 1.225 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 2.740 1.640 3.000 ;
        RECT  1.225 2.170 1.485 3.000 ;
        RECT  0.385 2.740 1.225 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX4MTH

MACRO INVX5MTH
    CLASS CORE ;
    FOREIGN INVX5MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 0.580 1.915 1.115 ;
        RECT  1.655 1.720 1.915 2.365 ;
        RECT  1.590 0.855 1.655 1.115 ;
        RECT  1.590 1.720 1.655 1.980 ;
        RECT  1.245 0.855 1.590 1.980 ;
        RECT  0.895 0.855 1.245 1.115 ;
        RECT  0.895 1.720 1.245 1.980 ;
        RECT  0.635 0.555 0.895 1.115 ;
        RECT  0.635 1.720 0.895 2.365 ;
        END
        AntennaDiffArea 0.966 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.295 1.065 1.540 ;
        END
        AntennaGateArea 0.5226 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 -0.130 2.050 0.130 ;
        RECT  1.145 -0.130 1.405 0.675 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.725 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 2.740 2.050 3.000 ;
        RECT  1.145 2.215 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.780 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX5MTH

MACRO INVX6MTH
    CLASS CORE ;
    FOREIGN INVX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 0.410 1.950 2.365 ;
        RECT  1.655 0.410 1.680 1.040 ;
        RECT  1.655 1.765 1.680 2.365 ;
        RECT  0.895 0.770 1.655 1.040 ;
        RECT  0.895 1.765 1.655 2.035 ;
        RECT  0.640 0.410 0.895 1.040 ;
        RECT  0.635 1.765 0.895 2.365 ;
        END
        AntennaDiffArea 1.137 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.290 1.485 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 -0.130 2.050 0.130 ;
        RECT  1.145 -0.130 1.405 0.590 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.405 2.740 2.050 3.000 ;
        RECT  1.145 2.215 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.780 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END INVX6MTH

MACRO INVX8MTH
    CLASS CORE ;
    FOREIGN INVX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 0.770 1.950 2.100 ;
        RECT  1.655 0.410 1.915 2.350 ;
        RECT  1.600 0.770 1.655 2.100 ;
        RECT  0.835 0.770 1.600 1.120 ;
        RECT  0.835 1.750 1.600 2.100 ;
        RECT  0.575 0.410 0.835 1.120 ;
        RECT  0.575 1.750 0.835 2.350 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.300 1.345 1.570 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.375 -0.130 2.460 0.130 ;
        RECT  1.115 -0.130 1.375 0.590 ;
        RECT  0.000 -0.130 1.115 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.375 2.740 2.460 3.000 ;
        RECT  1.115 2.280 1.375 3.000 ;
        RECT  0.000 2.740 1.115 3.000 ;
        END
    END VDD
END INVX8MTH

MACRO INVXLMTH
    CLASS CORE ;
    FOREIGN INVXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.765 1.130 2.035 ;
        RECT  0.710 0.765 0.920 1.025 ;
        RECT  0.680 1.760 0.920 2.035 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.210 0.720 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 -0.130 1.230 0.130 ;
        RECT  0.140 -0.130 0.400 1.025 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.400 2.740 1.230 3.000 ;
        RECT  0.140 1.825 0.400 3.000 ;
        RECT  0.000 2.740 0.140 3.000 ;
        END
    END VDD
END INVXLMTH

MACRO MDFFHQX1MTH
    CLASS CORE ;
    FOREIGN MDFFHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 1.025 2.435 1.540 ;
        END
        AntennaGateArea 0.1196 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.170 1.290 12.200 1.580 ;
        RECT  11.990 0.740 12.170 2.030 ;
        RECT  11.965 0.740 11.990 1.000 ;
        RECT  11.965 1.770 11.990 2.030 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 1.290 1.540 1.815 ;
        END
        AntennaGateArea 0.0611 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.485 0.470 3.590 0.770 ;
        RECT  3.325 0.470 3.485 1.250 ;
        RECT  3.295 0.990 3.325 1.250 ;
        END
        AntennaGateArea 0.0663 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.300 0.565 4.530 1.170 ;
        RECT  4.110 0.880 4.300 1.170 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.990 -0.130 12.300 0.130 ;
        RECT  11.610 -0.130 11.990 0.300 ;
        RECT  11.450 -0.130 11.610 0.965 ;
        RECT  11.390 -0.130 11.450 0.300 ;
        RECT  11.200 -0.130 11.390 0.130 ;
        RECT  10.260 -0.130 11.200 0.300 ;
        RECT  8.710 -0.130 10.260 0.130 ;
        RECT  8.110 -0.130 8.710 0.380 ;
        RECT  7.675 -0.130 8.110 0.130 ;
        RECT  7.415 -0.130 7.675 0.250 ;
        RECT  6.235 -0.130 7.415 0.130 ;
        RECT  5.735 -0.130 6.235 0.300 ;
        RECT  5.365 -0.130 5.735 0.130 ;
        RECT  4.425 -0.130 5.365 0.300 ;
        RECT  3.605 -0.130 4.425 0.130 ;
        RECT  3.005 -0.130 3.605 0.250 ;
        RECT  1.525 -0.130 3.005 0.130 ;
        RECT  1.265 -0.130 1.525 0.880 ;
        RECT  0.000 -0.130 1.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.635 2.740 12.300 3.000 ;
        RECT  11.035 2.400 11.635 3.000 ;
        RECT  10.835 2.740 11.035 3.000 ;
        RECT  10.305 2.395 10.835 3.000 ;
        RECT  3.205 2.740 10.305 3.000 ;
        RECT  2.705 2.570 3.205 3.000 ;
        RECT  0.000 2.740 2.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.110 0.600 11.270 2.110 ;
        RECT  10.880 0.600 11.110 0.760 ;
        RECT  10.995 1.575 11.110 2.110 ;
        RECT  10.535 1.575 10.995 1.735 ;
        RECT  10.730 0.940 10.890 1.235 ;
        RECT  10.000 0.940 10.730 1.100 ;
        RECT  10.375 1.460 10.535 1.735 ;
        RECT  10.005 2.270 10.105 2.430 ;
        RECT  9.845 2.060 10.005 2.430 ;
        RECT  9.840 0.545 10.000 1.855 ;
        RECT  9.465 2.060 9.845 2.220 ;
        RECT  9.565 0.545 9.840 0.705 ;
        RECT  9.645 1.695 9.840 1.855 ;
        RECT  9.465 0.920 9.655 1.145 ;
        RECT  6.750 2.400 9.485 2.560 ;
        RECT  9.395 0.920 9.465 2.220 ;
        RECT  9.305 0.985 9.395 2.220 ;
        RECT  9.215 0.545 9.315 0.705 ;
        RECT  7.090 2.060 9.305 2.220 ;
        RECT  9.125 0.545 9.215 0.760 ;
        RECT  9.055 0.545 9.125 1.860 ;
        RECT  8.965 0.600 9.055 1.860 ;
        RECT  8.305 0.600 8.965 0.760 ;
        RECT  8.865 1.700 8.965 1.860 ;
        RECT  8.685 1.030 8.785 1.290 ;
        RECT  8.525 1.030 8.685 1.810 ;
        RECT  7.965 1.650 8.525 1.810 ;
        RECT  8.145 0.600 8.305 1.265 ;
        RECT  7.805 0.650 7.965 1.810 ;
        RECT  7.435 0.650 7.805 0.810 ;
        RECT  7.435 1.650 7.805 1.810 ;
        RECT  7.090 1.010 7.615 1.270 ;
        RECT  7.275 0.550 7.435 0.810 ;
        RECT  7.275 1.620 7.435 1.880 ;
        RECT  6.930 0.600 7.090 2.220 ;
        RECT  6.055 0.600 6.930 0.760 ;
        RECT  6.590 1.000 6.750 2.560 ;
        RECT  6.260 1.000 6.590 1.160 ;
        RECT  6.060 1.960 6.590 2.120 ;
        RECT  6.250 2.300 6.410 2.560 ;
        RECT  3.545 2.400 6.250 2.560 ;
        RECT  5.900 1.960 6.060 2.220 ;
        RECT  5.895 0.600 6.055 1.745 ;
        RECT  3.885 2.060 5.900 2.220 ;
        RECT  5.425 0.600 5.895 0.760 ;
        RECT  5.775 1.280 5.895 1.745 ;
        RECT  5.445 1.585 5.775 1.745 ;
        RECT  4.965 1.170 5.555 1.330 ;
        RECT  5.175 1.585 5.445 1.850 ;
        RECT  4.965 0.590 5.175 0.850 ;
        RECT  4.550 1.690 5.175 1.850 ;
        RECT  4.805 0.590 4.965 1.510 ;
        RECT  4.370 1.350 4.805 1.510 ;
        RECT  4.210 1.350 4.370 1.835 ;
        RECT  4.065 1.575 4.210 1.835 ;
        RECT  3.930 0.540 4.115 0.700 ;
        RECT  3.885 0.540 3.930 1.355 ;
        RECT  3.770 0.540 3.885 2.220 ;
        RECT  3.725 1.145 3.770 2.220 ;
        RECT  3.385 2.110 3.545 2.560 ;
        RECT  2.775 2.110 3.385 2.270 ;
        RECT  3.115 0.610 3.145 0.890 ;
        RECT  2.955 0.610 3.115 1.930 ;
        RECT  2.095 0.310 2.805 0.470 ;
        RECT  2.615 0.680 2.775 2.270 ;
        RECT  2.345 0.680 2.615 0.840 ;
        RECT  2.525 1.720 2.615 2.270 ;
        RECT  2.365 1.720 2.525 2.560 ;
        RECT  0.335 2.400 2.365 2.560 ;
        RECT  1.920 1.905 2.140 2.220 ;
        RECT  1.935 0.310 2.095 0.800 ;
        RECT  1.920 0.640 1.935 0.800 ;
        RECT  1.760 0.640 1.920 2.220 ;
        RECT  0.675 2.060 1.760 2.220 ;
        RECT  0.855 0.640 1.015 1.880 ;
        RECT  0.695 0.640 0.855 0.800 ;
        RECT  0.515 1.250 0.675 2.220 ;
        RECT  0.445 1.250 0.515 1.510 ;
        RECT  0.265 0.590 0.335 0.850 ;
        RECT  0.265 1.880 0.335 2.560 ;
        RECT  0.105 0.590 0.265 2.560 ;
    END
END MDFFHQX1MTH

MACRO MDFFHQX2MTH
    CLASS CORE ;
    FOREIGN MDFFHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.070 1.025 2.360 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.555 1.290 12.610 1.580 ;
        RECT  12.375 0.425 12.555 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.220 1.125 1.540 1.580 ;
        RECT  1.195 1.125 1.220 1.385 ;
        END
        AntennaGateArea 0.0884 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.455 0.470 3.590 0.770 ;
        RECT  3.295 0.470 3.455 1.270 ;
        END
        AntennaGateArea 0.0871 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.260 0.680 4.530 1.170 ;
        RECT  4.110 0.920 4.260 1.170 ;
        END
        AntennaGateArea 0.1417 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.025 -0.130 12.710 0.130 ;
        RECT  11.865 -0.130 12.025 1.025 ;
        RECT  10.995 -0.130 11.865 0.130 ;
        RECT  10.395 -0.130 10.995 0.300 ;
        RECT  8.710 -0.130 10.395 0.130 ;
        RECT  7.770 -0.130 8.710 0.380 ;
        RECT  6.505 -0.130 7.770 0.130 ;
        RECT  5.565 -0.130 6.505 0.320 ;
        RECT  4.545 -0.130 5.565 0.130 ;
        RECT  4.285 -0.130 4.545 0.350 ;
        RECT  3.565 -0.130 4.285 0.130 ;
        RECT  3.305 -0.130 3.565 0.285 ;
        RECT  1.535 -0.130 3.305 0.130 ;
        RECT  1.275 -0.130 1.535 0.925 ;
        RECT  0.000 -0.130 1.275 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.025 2.740 12.710 3.000 ;
        RECT  11.865 1.775 12.025 3.000 ;
        RECT  11.685 2.740 11.865 3.000 ;
        RECT  10.745 2.435 11.685 3.000 ;
        RECT  3.205 2.740 10.745 3.000 ;
        RECT  2.705 2.570 3.205 3.000 ;
        RECT  0.000 2.740 2.705 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.460 0.565 11.620 2.145 ;
        RECT  11.305 0.565 11.460 0.725 ;
        RECT  11.355 1.725 11.460 2.145 ;
        RECT  10.845 1.725 11.355 1.885 ;
        RECT  11.110 1.010 11.270 1.290 ;
        RECT  10.375 1.130 11.110 1.290 ;
        RECT  10.585 1.560 10.845 1.885 ;
        RECT  10.215 0.595 10.375 1.875 ;
        RECT  10.265 2.365 10.365 2.525 ;
        RECT  10.105 2.060 10.265 2.525 ;
        RECT  10.130 0.595 10.215 0.755 ;
        RECT  9.680 1.715 10.215 1.875 ;
        RECT  9.530 0.495 10.130 0.755 ;
        RECT  9.495 2.060 10.105 2.220 ;
        RECT  9.760 0.935 10.020 1.195 ;
        RECT  6.755 2.400 9.885 2.560 ;
        RECT  9.495 1.035 9.760 1.195 ;
        RECT  9.335 1.035 9.495 2.220 ;
        RECT  7.095 2.060 9.335 2.220 ;
        RECT  9.150 0.580 9.250 0.840 ;
        RECT  8.990 0.580 9.150 1.875 ;
        RECT  8.330 0.680 8.990 0.840 ;
        RECT  8.855 1.715 8.990 1.875 ;
        RECT  8.675 1.120 8.810 1.380 ;
        RECT  8.515 1.120 8.675 1.610 ;
        RECT  7.990 1.450 8.515 1.610 ;
        RECT  8.170 0.680 8.330 1.265 ;
        RECT  7.830 0.650 7.990 1.610 ;
        RECT  7.435 0.650 7.830 0.810 ;
        RECT  7.435 1.450 7.830 1.610 ;
        RECT  7.095 1.010 7.635 1.270 ;
        RECT  7.275 0.550 7.435 0.810 ;
        RECT  7.275 1.450 7.435 1.880 ;
        RECT  6.935 0.630 7.095 2.220 ;
        RECT  6.055 0.630 6.935 0.790 ;
        RECT  6.595 1.000 6.755 2.560 ;
        RECT  6.445 1.000 6.595 1.160 ;
        RECT  6.060 1.960 6.595 2.120 ;
        RECT  6.255 2.300 6.415 2.560 ;
        RECT  3.545 2.400 6.255 2.560 ;
        RECT  6.055 1.310 6.155 1.470 ;
        RECT  5.900 1.960 6.060 2.220 ;
        RECT  5.895 0.630 6.055 1.745 ;
        RECT  3.885 2.060 5.900 2.220 ;
        RECT  5.365 0.630 5.895 0.790 ;
        RECT  5.445 1.585 5.895 1.745 ;
        RECT  4.875 1.170 5.555 1.330 ;
        RECT  5.175 1.585 5.445 1.850 ;
        RECT  4.600 1.690 5.175 1.850 ;
        RECT  4.875 0.580 5.115 0.740 ;
        RECT  4.715 0.580 4.875 1.510 ;
        RECT  4.370 1.350 4.715 1.510 ;
        RECT  4.210 1.350 4.370 1.830 ;
        RECT  4.065 1.570 4.210 1.830 ;
        RECT  3.930 0.580 4.075 0.740 ;
        RECT  3.885 0.580 3.930 1.355 ;
        RECT  3.770 0.580 3.885 2.220 ;
        RECT  3.725 1.145 3.770 2.220 ;
        RECT  3.385 2.230 3.545 2.560 ;
        RECT  2.700 2.230 3.385 2.390 ;
        RECT  3.115 1.640 3.205 1.900 ;
        RECT  2.955 0.630 3.115 1.900 ;
        RECT  2.925 1.640 2.955 1.900 ;
        RECT  2.145 0.310 2.825 0.470 ;
        RECT  2.540 0.680 2.700 2.390 ;
        RECT  2.395 0.680 2.540 0.840 ;
        RECT  2.525 1.760 2.540 2.390 ;
        RECT  2.365 1.760 2.525 2.560 ;
        RECT  0.335 2.400 2.365 2.560 ;
        RECT  1.885 1.760 2.185 2.220 ;
        RECT  1.985 0.310 2.145 0.825 ;
        RECT  1.885 0.665 1.985 0.825 ;
        RECT  1.725 0.665 1.885 2.220 ;
        RECT  0.675 2.060 1.725 2.220 ;
        RECT  1.015 1.620 1.040 1.880 ;
        RECT  0.855 0.710 1.015 1.880 ;
        RECT  0.730 0.710 0.855 0.870 ;
        RECT  0.515 1.325 0.675 2.220 ;
        RECT  0.485 1.325 0.515 1.585 ;
        RECT  0.305 0.665 0.430 0.925 ;
        RECT  0.305 1.720 0.335 2.560 ;
        RECT  0.145 0.665 0.305 2.560 ;
    END
END MDFFHQX2MTH

MACRO MDFFHQX4MTH
    CLASS CORE ;
    FOREIGN MDFFHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 1.085 2.360 1.580 ;
        RECT  1.880 1.085 2.085 1.245 ;
        RECT  1.720 0.430 1.880 1.245 ;
        RECT  0.680 0.430 1.720 0.590 ;
        RECT  0.520 0.430 0.680 1.245 ;
        END
        AntennaGateArea 0.2132 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.965 1.290 13.020 1.580 ;
        RECT  12.785 0.425 12.965 2.355 ;
        RECT  12.635 0.425 12.785 1.025 ;
        RECT  12.635 1.755 12.785 2.355 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.020 1.540 1.875 ;
        END
        AntennaGateArea 0.1599 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 0.470 4.000 0.760 ;
        RECT  3.705 0.470 3.865 1.250 ;
        END
        AntennaGateArea 0.1352 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.670 0.595 4.940 1.130 ;
        RECT  4.520 0.855 4.670 1.130 ;
        END
        AntennaGateArea 0.2015 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 -0.130 13.530 0.130 ;
        RECT  13.145 -0.130 13.405 1.025 ;
        RECT  12.355 -0.130 13.145 0.130 ;
        RECT  11.415 -0.130 12.355 0.300 ;
        RECT  11.200 -0.130 11.415 0.130 ;
        RECT  10.980 -0.130 11.200 0.855 ;
        RECT  10.495 -0.130 10.980 0.300 ;
        RECT  9.120 -0.130 10.495 0.130 ;
        RECT  8.860 -0.130 9.120 0.695 ;
        RECT  8.520 -0.130 8.860 0.345 ;
        RECT  6.810 -0.130 8.520 0.130 ;
        RECT  6.210 -0.130 6.810 0.375 ;
        RECT  2.370 -0.130 6.210 0.130 ;
        RECT  1.430 -0.130 2.370 0.250 ;
        RECT  0.000 -0.130 1.430 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.850 13.405 3.000 ;
        RECT  12.355 2.740 13.145 3.000 ;
        RECT  11.755 2.450 12.355 3.000 ;
        RECT  11.575 2.740 11.755 3.000 ;
        RECT  11.075 2.450 11.575 3.000 ;
        RECT  3.620 2.740 11.075 3.000 ;
        RECT  3.020 2.570 3.620 3.000 ;
        RECT  2.700 2.740 3.020 3.000 ;
        RECT  2.440 2.570 2.700 3.000 ;
        RECT  0.000 2.740 2.440 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.185 0.815 12.345 1.885 ;
        RECT  11.865 0.815 12.185 0.975 ;
        RECT  11.910 1.725 12.185 1.885 ;
        RECT  11.405 1.190 12.005 1.460 ;
        RECT  11.645 1.725 11.910 2.145 ;
        RECT  11.605 0.715 11.865 0.975 ;
        RECT  11.185 1.725 11.645 1.885 ;
        RECT  10.670 1.190 11.405 1.350 ;
        RECT  10.925 1.560 11.185 1.885 ;
        RECT  10.695 2.365 10.795 2.525 ;
        RECT  10.535 2.060 10.695 2.525 ;
        RECT  10.510 0.565 10.670 1.875 ;
        RECT  9.925 2.060 10.535 2.220 ;
        RECT  10.235 0.565 10.510 0.725 ;
        RECT  10.105 1.715 10.510 1.875 ;
        RECT  7.270 2.400 10.315 2.560 ;
        RECT  9.975 0.465 10.235 0.725 ;
        RECT  9.925 0.985 10.025 1.245 ;
        RECT  9.765 0.985 9.925 2.220 ;
        RECT  7.670 2.060 9.765 2.220 ;
        RECT  9.580 0.535 9.725 0.795 ;
        RECT  9.420 0.535 9.580 1.875 ;
        RECT  8.760 0.915 9.420 1.075 ;
        RECT  9.285 1.715 9.420 1.875 ;
        RECT  9.100 1.275 9.240 1.535 ;
        RECT  8.940 1.275 9.100 1.765 ;
        RECT  8.420 1.605 8.940 1.765 ;
        RECT  8.600 0.915 8.760 1.265 ;
        RECT  8.260 0.655 8.420 1.765 ;
        RECT  8.000 0.655 8.260 0.815 ;
        RECT  8.160 1.605 8.260 1.765 ;
        RECT  7.900 1.605 8.160 1.865 ;
        RECT  7.670 1.005 8.080 1.265 ;
        RECT  7.500 0.555 8.000 0.815 ;
        RECT  7.510 1.005 7.670 2.220 ;
        RECT  7.320 1.005 7.510 1.265 ;
        RECT  7.160 0.620 7.320 1.265 ;
        RECT  7.110 1.960 7.270 2.560 ;
        RECT  6.500 0.620 7.160 0.780 ;
        RECT  6.980 1.960 7.110 2.120 ;
        RECT  6.820 0.985 6.980 2.120 ;
        RECT  6.770 2.300 6.930 2.560 ;
        RECT  6.470 1.960 6.820 2.120 ;
        RECT  4.000 2.400 6.770 2.560 ;
        RECT  6.340 0.620 6.500 1.745 ;
        RECT  6.310 1.960 6.470 2.220 ;
        RECT  5.925 0.620 6.340 0.780 ;
        RECT  5.685 1.585 6.340 1.745 ;
        RECT  4.340 2.060 6.310 2.220 ;
        RECT  5.665 0.520 5.925 0.780 ;
        RECT  5.285 1.170 5.855 1.330 ;
        RECT  5.465 1.585 5.685 1.850 ;
        RECT  5.425 1.650 5.465 1.850 ;
        RECT  5.055 1.650 5.425 1.810 ;
        RECT  5.285 0.415 5.415 0.675 ;
        RECT  5.125 0.415 5.285 1.470 ;
        RECT  4.735 1.310 5.125 1.470 ;
        RECT  4.535 1.310 4.735 1.595 ;
        RECT  4.340 0.415 4.485 0.675 ;
        RECT  4.180 0.415 4.340 2.220 ;
        RECT  3.840 2.105 4.000 2.560 ;
        RECT  3.185 2.105 3.840 2.265 ;
        RECT  3.525 1.645 3.565 1.905 ;
        RECT  3.365 0.415 3.525 1.905 ;
        RECT  3.025 0.405 3.185 2.265 ;
        RECT  2.745 0.405 3.025 0.565 ;
        RECT  2.895 1.660 3.025 1.920 ;
        RECT  2.220 2.105 3.025 2.265 ;
        RECT  2.700 0.985 2.845 1.245 ;
        RECT  2.540 0.745 2.700 1.920 ;
        RECT  2.495 0.745 2.540 0.905 ;
        RECT  1.880 1.760 2.540 1.920 ;
        RECT  2.235 0.615 2.495 0.905 ;
        RECT  2.060 2.105 2.220 2.560 ;
        RECT  0.335 2.400 2.060 2.560 ;
        RECT  1.720 1.760 1.880 2.220 ;
        RECT  0.675 2.060 1.720 2.220 ;
        RECT  0.990 0.770 1.150 1.880 ;
        RECT  0.860 0.770 0.990 0.930 ;
        RECT  0.860 1.720 0.990 1.880 ;
        RECT  0.515 1.465 0.675 2.220 ;
        RECT  0.490 1.465 0.515 1.725 ;
        RECT  0.310 0.560 0.340 0.820 ;
        RECT  0.310 1.875 0.335 2.560 ;
        RECT  0.150 0.560 0.310 2.560 ;
    END
END MDFFHQX4MTH

MACRO MDFFHQX8MTH
    CLASS CORE ;
    FOREIGN MDFFHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.130 2.230 1.580 ;
        RECT  1.740 0.770 1.900 1.580 ;
        RECT  1.455 0.770 1.740 0.930 ;
        RECT  1.295 0.325 1.455 0.930 ;
        RECT  0.675 0.325 1.295 0.485 ;
        RECT  0.515 0.325 0.675 1.245 ;
        END
        AntennaGateArea 0.2132 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.755 1.685 13.825 2.285 ;
        RECT  13.495 0.425 13.755 2.285 ;
        RECT  12.755 1.290 13.495 1.580 ;
        RECT  12.735 1.290 12.755 2.285 ;
        RECT  12.475 0.425 12.735 2.285 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.160 1.545 1.875 ;
        END
        AntennaGateArea 0.1599 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 0.470 4.000 0.760 ;
        RECT  3.705 0.470 3.865 1.250 ;
        END
        AntennaGateArea 0.1352 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.670 0.595 4.940 1.130 ;
        RECT  4.520 0.880 4.670 1.130 ;
        END
        AntennaGateArea 0.2015 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.175 -0.130 14.350 0.130 ;
        RECT  13.975 -0.130 14.175 1.025 ;
        RECT  13.175 -0.130 13.975 0.130 ;
        RECT  12.955 -0.130 13.175 1.025 ;
        RECT  12.095 -0.130 12.955 0.130 ;
        RECT  11.595 -0.130 12.095 0.300 ;
        RECT  11.150 -0.130 11.595 0.130 ;
        RECT  10.930 -0.130 11.150 0.855 ;
        RECT  10.495 -0.130 10.930 0.300 ;
        RECT  9.120 -0.130 10.495 0.130 ;
        RECT  8.520 -0.130 9.120 0.300 ;
        RECT  6.755 -0.130 8.520 0.130 ;
        RECT  6.255 -0.130 6.755 0.300 ;
        RECT  2.250 -0.130 6.255 0.130 ;
        RECT  1.910 -0.130 2.250 0.360 ;
        RECT  1.650 -0.130 1.910 0.545 ;
        RECT  0.000 -0.130 1.650 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.295 2.740 14.350 3.000 ;
        RECT  13.075 1.770 13.295 3.000 ;
        RECT  12.265 2.740 13.075 3.000 ;
        RECT  11.660 2.450 12.265 3.000 ;
        RECT  11.475 2.740 11.660 3.000 ;
        RECT  11.210 2.450 11.475 3.000 ;
        RECT  3.540 2.740 11.210 3.000 ;
        RECT  2.940 2.570 3.540 3.000 ;
        RECT  2.720 2.740 2.940 3.000 ;
        RECT  2.460 2.565 2.720 3.000 ;
        RECT  0.000 2.740 2.460 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.070 0.805 12.230 1.885 ;
        RECT  11.770 0.805 12.070 0.965 ;
        RECT  11.900 1.725 12.070 1.885 ;
        RECT  11.685 1.725 11.900 2.145 ;
        RECT  11.390 1.190 11.890 1.450 ;
        RECT  11.510 0.705 11.770 0.965 ;
        RECT  11.055 1.725 11.685 1.885 ;
        RECT  10.670 1.190 11.390 1.350 ;
        RECT  10.895 1.560 11.055 1.885 ;
        RECT  10.695 2.365 10.795 2.525 ;
        RECT  10.535 2.060 10.695 2.525 ;
        RECT  10.510 0.565 10.670 1.875 ;
        RECT  9.925 2.060 10.535 2.220 ;
        RECT  10.235 0.565 10.510 0.725 ;
        RECT  10.105 1.715 10.510 1.875 ;
        RECT  7.345 2.400 10.315 2.560 ;
        RECT  9.975 0.465 10.235 0.725 ;
        RECT  9.925 1.035 10.025 1.195 ;
        RECT  9.765 1.035 9.925 2.220 ;
        RECT  7.685 2.060 9.765 2.220 ;
        RECT  9.580 0.580 9.725 0.840 ;
        RECT  9.465 0.580 9.580 1.875 ;
        RECT  9.420 0.680 9.465 1.875 ;
        RECT  8.760 0.680 9.420 0.840 ;
        RECT  9.285 1.715 9.420 1.875 ;
        RECT  9.100 1.190 9.240 1.450 ;
        RECT  8.940 1.190 9.100 1.765 ;
        RECT  8.420 1.605 8.940 1.765 ;
        RECT  8.600 0.680 8.760 1.265 ;
        RECT  8.260 0.655 8.420 1.765 ;
        RECT  8.080 0.655 8.260 0.815 ;
        RECT  8.110 1.605 8.260 1.765 ;
        RECT  7.950 1.605 8.110 1.865 ;
        RECT  7.920 0.555 8.080 0.815 ;
        RECT  7.685 1.005 8.080 1.265 ;
        RECT  7.525 0.620 7.685 2.220 ;
        RECT  6.525 0.620 7.525 0.780 ;
        RECT  7.185 1.035 7.345 2.560 ;
        RECT  6.865 1.035 7.185 1.195 ;
        RECT  6.470 1.960 7.185 2.120 ;
        RECT  3.930 2.400 7.005 2.560 ;
        RECT  6.365 0.620 6.525 1.745 ;
        RECT  6.310 1.960 6.470 2.220 ;
        RECT  5.925 0.620 6.365 0.780 ;
        RECT  5.795 1.585 6.365 1.745 ;
        RECT  4.340 2.060 6.310 2.220 ;
        RECT  5.285 1.170 5.965 1.330 ;
        RECT  5.665 0.520 5.925 0.780 ;
        RECT  5.535 1.585 5.795 1.880 ;
        RECT  5.165 1.720 5.535 1.880 ;
        RECT  5.285 0.465 5.415 0.625 ;
        RECT  5.125 0.465 5.285 1.495 ;
        RECT  4.735 1.335 5.125 1.495 ;
        RECT  4.535 1.335 4.735 1.595 ;
        RECT  4.340 0.415 4.435 0.675 ;
        RECT  4.180 0.415 4.340 2.220 ;
        RECT  3.770 2.105 3.930 2.560 ;
        RECT  3.185 2.105 3.770 2.265 ;
        RECT  3.525 1.645 3.565 1.905 ;
        RECT  3.365 0.415 3.525 1.905 ;
        RECT  3.025 0.405 3.185 2.265 ;
        RECT  2.730 0.405 3.025 0.565 ;
        RECT  2.895 1.660 3.025 2.265 ;
        RECT  2.250 2.105 2.895 2.265 ;
        RECT  2.685 0.985 2.830 1.245 ;
        RECT  2.525 0.740 2.685 1.920 ;
        RECT  2.430 0.740 2.525 0.900 ;
        RECT  1.885 1.760 2.525 1.920 ;
        RECT  2.270 0.615 2.430 0.900 ;
        RECT  2.090 2.105 2.250 2.560 ;
        RECT  0.335 2.400 2.090 2.560 ;
        RECT  1.725 1.760 1.885 2.220 ;
        RECT  0.675 2.060 1.725 2.220 ;
        RECT  1.015 0.665 1.115 0.825 ;
        RECT  1.015 1.620 1.055 1.880 ;
        RECT  0.855 0.665 1.015 1.880 ;
        RECT  0.515 1.465 0.675 2.220 ;
        RECT  0.475 1.465 0.515 1.725 ;
        RECT  0.295 0.560 0.335 0.820 ;
        RECT  0.295 1.995 0.335 2.560 ;
        RECT  0.135 0.560 0.295 2.560 ;
    END
END MDFFHQX8MTH

MACRO MX2X12MTH
    CLASS CORE ;
    FOREIGN MX2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.075 0.405 6.335 2.290 ;
        RECT  5.315 1.065 6.075 1.785 ;
        RECT  5.055 0.405 5.315 2.290 ;
        RECT  4.305 0.465 5.055 1.005 ;
        RECT  4.355 1.690 5.055 2.230 ;
        RECT  4.145 1.690 4.355 2.290 ;
        RECT  4.145 0.405 4.305 1.005 ;
        END
        AntennaDiffArea 1.8 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 1.315 2.745 2.125 ;
        RECT  2.245 1.965 2.585 2.125 ;
        RECT  2.085 1.965 2.245 2.435 ;
        RECT  1.755 2.275 2.085 2.435 ;
        RECT  1.495 2.275 1.755 2.540 ;
        RECT  0.555 2.275 1.495 2.435 ;
        RECT  0.100 2.110 0.555 2.435 ;
        END
        AntennaGateArea 0.2925 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.850 0.880 1.130 1.405 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.110 3.285 1.650 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 -0.130 6.970 0.130 ;
        RECT  6.585 -0.130 6.845 0.945 ;
        RECT  5.825 -0.130 6.585 0.130 ;
        RECT  5.565 -0.130 5.825 0.835 ;
        RECT  3.815 -0.130 5.565 0.130 ;
        RECT  3.215 -0.130 3.815 0.250 ;
        RECT  0.915 -0.130 3.215 0.130 ;
        RECT  0.315 -0.130 0.915 0.350 ;
        RECT  0.000 -0.130 0.315 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 1.965 6.845 3.000 ;
        RECT  5.825 2.740 6.585 3.000 ;
        RECT  5.565 1.965 5.825 3.000 ;
        RECT  3.755 2.740 5.565 3.000 ;
        RECT  3.495 2.535 3.755 3.000 ;
        RECT  0.845 2.740 3.495 3.000 ;
        RECT  0.245 2.615 0.845 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.965 1.185 4.865 1.345 ;
        RECT  3.805 0.430 3.965 2.355 ;
        RECT  2.065 0.430 3.805 0.590 ;
        RECT  3.280 2.195 3.805 2.355 ;
        RECT  3.465 0.770 3.625 2.015 ;
        RECT  2.640 0.770 3.465 0.930 ;
        RECT  2.935 1.855 3.465 2.015 ;
        RECT  3.030 2.195 3.280 2.490 ;
        RECT  2.685 2.330 3.030 2.490 ;
        RECT  2.425 2.305 2.685 2.490 ;
        RECT  2.245 0.845 2.405 1.785 ;
        RECT  1.470 0.845 2.245 1.005 ;
        RECT  1.905 1.625 2.245 1.785 ;
        RECT  1.805 0.380 2.065 0.640 ;
        RECT  1.905 1.185 2.065 1.445 ;
        RECT  1.565 1.285 1.905 1.445 ;
        RECT  1.745 1.625 1.905 2.090 ;
        RECT  1.125 1.930 1.745 2.090 ;
        RECT  1.405 1.285 1.565 1.750 ;
        RECT  1.310 0.440 1.470 1.005 ;
        RECT  0.385 1.590 1.405 1.750 ;
        RECT  1.195 0.440 1.310 0.700 ;
        RECT  0.285 0.765 0.385 1.025 ;
        RECT  0.285 1.590 0.385 1.920 ;
        RECT  0.125 0.765 0.285 1.920 ;
    END
END MX2X12MTH

MACRO MX2X1MTH
    CLASS CORE ;
    FOREIGN MX2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.765 0.550 4.000 2.285 ;
        END
        AntennaDiffArea 0.34 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.400 1.580 ;
        END
        AntennaGateArea 0.1612 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.280 1.435 ;
        END
        AntennaGateArea 0.1079 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 1.290 3.245 1.675 ;
        END
        AntennaGateArea 0.1079 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.415 -0.130 4.100 0.130 ;
        RECT  3.255 -0.130 3.415 0.770 ;
        RECT  3.155 -0.130 3.255 0.250 ;
        RECT  1.155 -0.130 3.155 0.130 ;
        RECT  0.895 -0.130 1.155 0.700 ;
        RECT  0.585 -0.130 0.895 0.130 ;
        RECT  0.325 -0.130 0.585 0.250 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.400 2.740 4.100 3.000 ;
        RECT  2.795 2.535 3.400 3.000 ;
        RECT  1.215 2.740 2.795 3.000 ;
        RECT  0.955 1.955 1.215 3.000 ;
        RECT  0.615 2.740 0.955 3.000 ;
        RECT  0.355 2.620 0.615 3.000 ;
        RECT  0.000 2.740 0.355 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.425 0.950 3.585 2.355 ;
        RECT  3.075 0.950 3.425 1.110 ;
        RECT  2.555 2.195 3.425 2.355 ;
        RECT  2.915 0.420 3.075 1.110 ;
        RECT  2.245 0.420 2.915 0.580 ;
        RECT  2.640 1.855 2.830 2.015 ;
        RECT  2.640 0.760 2.735 1.020 ;
        RECT  2.480 0.760 2.640 2.015 ;
        RECT  2.395 2.195 2.555 2.455 ;
        RECT  2.030 2.295 2.395 2.455 ;
        RECT  1.985 0.420 2.245 0.795 ;
        RECT  2.055 0.975 2.215 2.115 ;
        RECT  1.725 0.975 2.055 1.135 ;
        RECT  1.480 1.955 2.055 2.115 ;
        RECT  1.710 1.315 1.870 1.775 ;
        RECT  1.465 0.645 1.725 1.135 ;
        RECT  0.740 1.615 1.710 1.775 ;
        RECT  0.615 0.815 0.740 1.955 ;
        RECT  0.580 0.815 0.615 2.055 ;
        RECT  0.320 0.715 0.580 0.975 ;
        RECT  0.355 1.795 0.580 2.055 ;
    END
END MX2X1MTH

MACRO MX2X2MTH
    CLASS CORE ;
    FOREIGN MX2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.765 0.405 4.000 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.400 1.580 ;
        END
        AntennaGateArea 0.247 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 1.205 1.495 1.435 ;
        RECT  0.920 0.880 1.210 1.435 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.820 1.290 3.245 1.675 ;
        END
        AntennaGateArea 0.1755 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 -0.130 4.100 0.130 ;
        RECT  3.255 -0.130 3.435 0.770 ;
        RECT  3.175 -0.130 3.255 0.250 ;
        RECT  1.185 -0.130 3.175 0.130 ;
        RECT  0.925 -0.130 1.185 0.700 ;
        RECT  0.615 -0.130 0.925 0.130 ;
        RECT  0.355 -0.130 0.615 0.250 ;
        RECT  0.000 -0.130 0.355 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  3.170 2.535 3.435 3.000 ;
        RECT  1.320 2.740 3.170 3.000 ;
        RECT  0.920 2.005 1.320 3.000 ;
        RECT  0.720 2.140 0.920 3.000 ;
        RECT  0.410 2.740 0.720 3.000 ;
        RECT  0.150 2.620 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.425 0.950 3.585 2.355 ;
        RECT  3.075 0.950 3.425 1.110 ;
        RECT  2.975 2.195 3.425 2.355 ;
        RECT  2.915 0.410 3.075 1.110 ;
        RECT  2.815 2.195 2.975 2.455 ;
        RECT  2.245 0.410 2.915 0.570 ;
        RECT  2.640 1.855 2.890 2.015 ;
        RECT  2.120 2.295 2.815 2.455 ;
        RECT  2.640 0.750 2.735 1.010 ;
        RECT  2.480 0.750 2.640 2.015 ;
        RECT  2.140 0.855 2.300 2.115 ;
        RECT  1.985 0.410 2.245 0.675 ;
        RECT  1.725 0.855 2.140 1.015 ;
        RECT  1.570 1.955 2.140 2.115 ;
        RECT  1.800 1.315 1.960 1.775 ;
        RECT  0.740 1.615 1.800 1.775 ;
        RECT  1.465 0.645 1.725 1.015 ;
        RECT  0.580 0.815 0.740 1.945 ;
        RECT  0.350 0.815 0.580 0.975 ;
        RECT  0.180 1.785 0.580 1.945 ;
    END
END MX2X2MTH

MACRO MX2X3MTH
    CLASS CORE ;
    FOREIGN MX2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 0.915 4.410 1.940 ;
        RECT  3.935 0.915 4.200 1.075 ;
        RECT  3.985 1.780 4.200 1.940 ;
        RECT  3.725 1.780 3.985 2.120 ;
        RECT  3.720 0.660 3.935 1.075 ;
        END
        AntennaDiffArea 0.472 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.645 2.380 1.745 2.540 ;
        RECT  1.485 2.195 1.645 2.540 ;
        RECT  0.555 2.195 1.485 2.355 ;
        RECT  0.100 2.110 0.555 2.400 ;
        END
        AntennaGateArea 0.286 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.715 0.880 1.135 1.305 ;
        END
        AntennaGateArea 0.2002 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.110 3.180 1.675 ;
        END
        AntennaGateArea 0.2002 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  4.125 -0.130 4.385 0.310 ;
        RECT  3.390 -0.130 4.125 0.130 ;
        RECT  3.130 -0.130 3.390 0.250 ;
        RECT  0.885 -0.130 3.130 0.130 ;
        RECT  0.285 -0.130 0.885 0.435 ;
        RECT  0.000 -0.130 0.285 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 2.570 4.385 3.000 ;
        RECT  0.835 2.740 4.125 3.000 ;
        RECT  0.235 2.585 0.835 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.520 1.255 4.020 1.515 ;
        RECT  3.360 0.430 3.520 2.355 ;
        RECT  1.685 0.430 3.360 0.590 ;
        RECT  2.495 2.195 3.360 2.355 ;
        RECT  2.715 1.855 3.005 2.015 ;
        RECT  2.715 0.770 2.815 0.930 ;
        RECT  2.555 0.770 2.715 2.015 ;
        RECT  2.235 2.195 2.495 2.455 ;
        RECT  2.215 0.770 2.375 2.015 ;
        RECT  1.475 0.770 2.215 0.930 ;
        RECT  1.115 1.855 2.215 2.015 ;
        RECT  1.875 1.110 2.035 1.370 ;
        RECT  1.475 1.210 1.875 1.370 ;
        RECT  1.315 0.400 1.475 0.930 ;
        RECT  1.315 1.210 1.475 1.645 ;
        RECT  1.165 0.400 1.315 0.660 ;
        RECT  0.385 1.485 1.315 1.645 ;
        RECT  0.225 0.725 0.385 1.930 ;
        RECT  0.125 0.725 0.225 0.985 ;
        RECT  0.125 1.770 0.225 1.930 ;
    END
END MX2X3MTH

MACRO MX2X4MTH
    CLASS CORE ;
    FOREIGN MX2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 1.290 4.410 1.580 ;
        RECT  4.180 0.840 4.285 1.710 ;
        RECT  4.105 0.840 4.180 2.290 ;
        RECT  4.090 0.840 4.105 1.000 ;
        RECT  3.965 1.525 4.105 2.290 ;
        RECT  3.875 0.400 4.090 1.000 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 2.275 1.835 2.540 ;
        RECT  0.505 2.275 1.575 2.435 ;
        RECT  0.100 2.110 0.505 2.435 ;
        END
        AntennaGateArea 0.286 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 0.880 1.130 1.405 ;
        END
        AntennaGateArea 0.2002 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.200 3.295 1.670 ;
        END
        AntennaGateArea 0.2002 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 -0.130 4.920 0.130 ;
        RECT  4.465 -0.130 4.725 0.905 ;
        RECT  3.545 -0.130 4.465 0.130 ;
        RECT  3.285 -0.130 3.545 0.250 ;
        RECT  0.925 -0.130 3.285 0.130 ;
        RECT  0.665 -0.130 0.925 0.595 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.715 2.740 4.920 3.000 ;
        RECT  4.455 1.890 4.715 3.000 ;
        RECT  3.635 2.740 4.455 3.000 ;
        RECT  3.375 2.535 3.635 3.000 ;
        RECT  0.945 2.740 3.375 3.000 ;
        RECT  0.325 2.615 0.945 3.000 ;
        RECT  0.000 2.740 0.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.695 1.185 3.915 1.345 ;
        RECT  3.535 0.430 3.695 2.355 ;
        RECT  2.445 0.430 3.535 0.590 ;
        RECT  2.325 2.195 3.535 2.355 ;
        RECT  2.790 1.855 3.095 2.015 ;
        RECT  2.790 0.770 2.955 0.930 ;
        RECT  2.630 0.770 2.790 2.015 ;
        RECT  2.290 0.855 2.450 1.975 ;
        RECT  1.845 0.430 2.445 0.675 ;
        RECT  1.500 0.855 2.290 1.015 ;
        RECT  2.035 1.815 2.290 1.975 ;
        RECT  1.950 1.195 2.110 1.635 ;
        RECT  1.815 1.815 2.035 2.090 ;
        RECT  1.505 1.475 1.950 1.635 ;
        RECT  1.205 1.930 1.815 2.090 ;
        RECT  1.310 1.475 1.505 1.750 ;
        RECT  1.340 0.380 1.500 1.015 ;
        RECT  1.235 0.380 1.340 0.640 ;
        RECT  0.685 1.590 1.310 1.750 ;
        RECT  0.525 0.775 0.685 1.920 ;
        RECT  0.125 0.775 0.525 0.935 ;
        RECT  0.125 1.760 0.525 1.920 ;
    END
END MX2X4MTH

MACRO MX2X6MTH
    CLASS CORE ;
    FOREIGN MX2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.195 0.845 5.230 1.785 ;
        RECT  4.935 0.405 5.195 2.290 ;
        RECT  4.115 0.775 4.935 1.005 ;
        RECT  4.180 1.525 4.935 1.785 ;
        RECT  3.915 1.525 4.180 2.290 ;
        RECT  3.855 0.405 4.115 1.005 ;
        END
        AntennaDiffArea 1.137 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.575 2.275 1.835 2.540 ;
        RECT  0.555 2.275 1.575 2.435 ;
        RECT  0.355 2.175 0.555 2.435 ;
        RECT  0.100 2.110 0.355 2.435 ;
        END
        AntennaGateArea 0.286 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 0.880 1.135 1.405 ;
        END
        AntennaGateArea 0.2002 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.110 3.335 1.670 ;
        END
        AntennaGateArea 0.2002 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.655 -0.130 5.330 0.130 ;
        RECT  4.395 -0.130 4.655 0.590 ;
        RECT  3.500 -0.130 4.395 0.130 ;
        RECT  3.240 -0.130 3.500 0.250 ;
        RECT  0.925 -0.130 3.240 0.130 ;
        RECT  0.665 -0.130 0.925 0.645 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.685 2.740 5.330 3.000 ;
        RECT  4.425 1.965 4.685 3.000 ;
        RECT  3.635 2.740 4.425 3.000 ;
        RECT  3.375 2.535 3.635 3.000 ;
        RECT  0.925 2.740 3.375 3.000 ;
        RECT  0.325 2.615 0.925 3.000 ;
        RECT  0.000 2.740 0.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.675 1.185 4.685 1.345 ;
        RECT  3.515 0.430 3.675 2.355 ;
        RECT  2.360 0.430 3.515 0.590 ;
        RECT  2.325 2.195 3.515 2.355 ;
        RECT  2.790 1.855 3.095 2.015 ;
        RECT  2.790 0.770 2.890 0.930 ;
        RECT  2.630 0.770 2.790 2.015 ;
        RECT  2.290 0.855 2.450 1.975 ;
        RECT  1.760 0.430 2.360 0.675 ;
        RECT  1.500 0.855 2.290 1.015 ;
        RECT  2.035 1.815 2.290 1.975 ;
        RECT  1.950 1.195 2.110 1.635 ;
        RECT  1.775 1.815 2.035 2.090 ;
        RECT  1.505 1.475 1.950 1.635 ;
        RECT  1.205 1.930 1.775 2.090 ;
        RECT  1.310 1.475 1.505 1.750 ;
        RECT  1.340 0.440 1.500 1.015 ;
        RECT  1.235 0.440 1.340 0.700 ;
        RECT  0.690 1.590 1.310 1.750 ;
        RECT  0.530 0.825 0.690 1.920 ;
        RECT  0.385 0.825 0.530 0.985 ;
        RECT  0.125 1.760 0.530 1.920 ;
        RECT  0.125 0.725 0.385 0.985 ;
    END
END MX2X6MTH

MACRO MX2X8MTH
    CLASS CORE ;
    FOREIGN MX2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.085 5.230 1.785 ;
        RECT  5.105 0.745 5.150 1.785 ;
        RECT  4.845 0.405 5.105 2.355 ;
        RECT  4.775 0.745 4.845 1.785 ;
        RECT  4.090 0.745 4.775 1.005 ;
        RECT  4.090 1.525 4.775 1.785 ;
        RECT  3.825 0.405 4.090 1.005 ;
        RECT  3.825 1.525 4.090 2.305 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 2.275 1.745 2.540 ;
        RECT  0.555 2.275 1.485 2.435 ;
        RECT  0.355 2.175 0.555 2.435 ;
        RECT  0.100 2.110 0.355 2.435 ;
        END
        AntennaGateArea 0.286 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 0.880 1.135 1.405 ;
        END
        AntennaGateArea 0.2002 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.110 3.295 1.670 ;
        END
        AntennaGateArea 0.2002 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 0.905 ;
        RECT  4.595 -0.130 5.355 0.130 ;
        RECT  4.335 -0.130 4.595 0.565 ;
        RECT  3.505 -0.130 4.335 0.130 ;
        RECT  3.245 -0.130 3.505 0.250 ;
        RECT  0.925 -0.130 3.245 0.130 ;
        RECT  0.665 -0.130 0.925 0.645 ;
        RECT  0.325 -0.130 0.665 0.305 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 1.965 5.615 3.000 ;
        RECT  4.595 2.740 5.355 3.000 ;
        RECT  4.335 1.965 4.595 3.000 ;
        RECT  3.545 2.740 4.335 3.000 ;
        RECT  3.285 2.535 3.545 3.000 ;
        RECT  0.855 2.740 3.285 3.000 ;
        RECT  0.235 2.615 0.855 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.645 1.185 4.595 1.345 ;
        RECT  3.485 0.430 3.645 2.355 ;
        RECT  2.360 0.430 3.485 0.590 ;
        RECT  2.235 2.195 3.485 2.355 ;
        RECT  2.790 1.855 3.005 2.015 ;
        RECT  2.790 0.770 2.890 0.930 ;
        RECT  2.630 0.770 2.790 2.015 ;
        RECT  2.290 0.855 2.450 1.975 ;
        RECT  1.760 0.430 2.360 0.675 ;
        RECT  1.500 0.855 2.290 1.015 ;
        RECT  1.945 1.815 2.290 1.975 ;
        RECT  1.950 1.195 2.110 1.635 ;
        RECT  1.505 1.475 1.950 1.635 ;
        RECT  1.685 1.815 1.945 2.090 ;
        RECT  1.115 1.930 1.685 2.090 ;
        RECT  1.310 1.475 1.505 1.750 ;
        RECT  1.340 0.440 1.500 1.015 ;
        RECT  1.240 0.440 1.340 0.700 ;
        RECT  0.695 1.590 1.310 1.750 ;
        RECT  0.535 0.825 0.695 1.920 ;
        RECT  0.385 0.825 0.535 0.985 ;
        RECT  0.125 1.760 0.535 1.920 ;
        RECT  0.125 0.725 0.385 0.985 ;
    END
END MX2X8MTH

MACRO MX2XLMTH
    CLASS CORE ;
    FOREIGN MX2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.765 4.000 2.145 ;
        RECT  3.715 0.765 3.790 1.025 ;
        RECT  3.735 1.885 3.790 2.145 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.865 1.500 2.025 1.760 ;
        RECT  1.465 1.500 1.865 1.660 ;
        RECT  1.305 0.695 1.465 1.660 ;
        RECT  0.565 0.920 1.305 1.130 ;
        RECT  0.465 0.970 0.565 1.130 ;
        END
        AntennaGateArea 0.1131 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.330 1.015 1.680 ;
        END
        AntennaGateArea 0.0598 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 1.290 2.855 1.755 ;
        END
        AntennaGateArea 0.0598 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 -0.130 4.100 0.130 ;
        RECT  3.280 -0.130 3.880 0.250 ;
        RECT  3.100 -0.130 3.280 0.130 ;
        RECT  2.500 -0.130 3.100 0.250 ;
        RECT  0.815 -0.130 2.500 0.130 ;
        RECT  0.555 -0.130 0.815 0.300 ;
        RECT  0.000 -0.130 0.555 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.935 2.740 4.100 3.000 ;
        RECT  3.335 2.620 3.935 3.000 ;
        RECT  3.155 2.740 3.335 3.000 ;
        RECT  2.215 2.620 3.155 3.000 ;
        RECT  1.205 2.740 2.215 3.000 ;
        RECT  0.265 2.620 1.205 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.535 1.185 3.610 1.445 ;
        RECT  3.375 0.475 3.535 2.440 ;
        RECT  2.145 0.475 3.375 0.635 ;
        RECT  1.915 2.280 3.375 2.440 ;
        RECT  3.035 0.815 3.195 2.095 ;
        RECT  2.505 0.815 3.035 0.975 ;
        RECT  2.545 1.935 3.035 2.095 ;
        RECT  2.205 1.160 2.365 2.100 ;
        RECT  1.805 1.160 2.205 1.320 ;
        RECT  1.125 1.940 2.205 2.100 ;
        RECT  1.985 0.475 2.145 0.980 ;
        RECT  1.755 2.280 1.915 2.540 ;
        RECT  1.645 0.355 1.805 1.320 ;
        RECT  1.145 0.355 1.645 0.515 ;
        RECT  1.385 2.280 1.545 2.560 ;
        RECT  0.385 2.280 1.385 2.440 ;
        RECT  0.285 0.530 0.385 0.790 ;
        RECT  0.285 1.885 0.385 2.440 ;
        RECT  0.225 0.530 0.285 2.440 ;
        RECT  0.125 0.530 0.225 2.145 ;
    END
END MX2XLMTH

MACRO MX3X1MTH
    CLASS CORE ;
    FOREIGN MX3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 1.290 6.050 1.580 ;
        RECT  5.825 0.805 6.025 2.085 ;
        RECT  5.765 0.805 5.825 1.005 ;
        RECT  5.765 1.825 5.825 2.085 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 1.075 3.255 1.530 ;
        RECT  2.970 1.075 3.180 1.580 ;
        END
        AntennaGateArea 0.1911 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.075 0.515 2.510 ;
        END
        AntennaGateArea 0.2184 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.325 1.290 5.640 1.580 ;
        RECT  5.165 1.145 5.325 1.580 ;
        END
        AntennaGateArea 0.1079 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.740 0.920 1.065 1.345 ;
        RECT  0.470 0.920 0.740 1.130 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 1.075 2.790 1.580 ;
        RECT  2.455 1.255 2.570 1.580 ;
        END
        AntennaGateArea 0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.485 -0.130 6.150 0.130 ;
        RECT  4.885 -0.130 5.485 0.250 ;
        RECT  0.955 -0.130 4.885 0.130 ;
        RECT  0.695 -0.130 0.955 0.740 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.485 2.740 6.150 3.000 ;
        RECT  4.885 2.455 5.485 3.000 ;
        RECT  3.445 2.740 4.885 3.000 ;
        RECT  2.845 2.550 3.445 3.000 ;
        RECT  0.955 2.740 2.845 3.000 ;
        RECT  0.695 1.945 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.665 0.375 5.925 0.590 ;
        RECT  4.535 0.430 5.665 0.590 ;
        RECT  4.955 0.770 5.065 0.930 ;
        RECT  4.955 1.915 5.065 2.075 ;
        RECT  4.795 0.770 4.955 2.075 ;
        RECT  4.375 0.430 4.535 2.145 ;
        RECT  4.345 0.720 4.375 0.980 ;
        RECT  4.345 1.885 4.375 2.145 ;
        RECT  3.995 0.665 4.045 1.605 ;
        RECT  3.945 0.665 3.995 2.365 ;
        RECT  3.885 0.395 3.945 2.365 ;
        RECT  3.785 0.395 3.885 0.865 ;
        RECT  3.835 1.445 3.885 2.365 ;
        RECT  1.755 2.205 3.835 2.365 ;
        RECT  2.045 0.395 3.785 0.555 ;
        RECT  3.595 1.105 3.695 1.265 ;
        RECT  3.435 0.735 3.595 1.995 ;
        RECT  3.275 0.735 3.435 0.895 ;
        RECT  3.325 1.735 3.435 1.995 ;
        RECT  2.385 0.735 2.555 0.895 ;
        RECT  2.345 1.760 2.505 2.020 ;
        RECT  2.275 0.735 2.385 1.075 ;
        RECT  2.275 1.760 2.345 1.920 ;
        RECT  2.225 0.735 2.275 1.920 ;
        RECT  2.115 0.915 2.225 1.920 ;
        RECT  1.885 0.395 2.045 0.735 ;
        RECT  1.775 0.975 1.935 2.025 ;
        RECT  1.785 0.575 1.885 0.735 ;
        RECT  1.455 0.975 1.775 1.135 ;
        RECT  1.215 1.865 1.775 2.025 ;
        RECT  1.435 1.315 1.595 1.685 ;
        RECT  1.295 0.655 1.455 1.135 ;
        RECT  0.385 1.525 1.435 1.685 ;
        RECT  0.285 0.580 0.385 0.740 ;
        RECT  0.285 1.525 0.385 1.895 ;
        RECT  0.125 0.580 0.285 1.895 ;
    END
END MX3X1MTH

MACRO MX3X2MTH
    CLASS CORE ;
    FOREIGN MX3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 0.485 7.280 2.495 ;
        RECT  6.995 1.895 7.045 2.495 ;
        END
        AntennaDiffArea 0.493 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.675 1.115 5.730 1.375 ;
        RECT  5.515 1.115 5.675 2.215 ;
        RECT  4.485 2.055 5.515 2.215 ;
        RECT  4.325 2.055 4.485 2.365 ;
        RECT  3.815 2.095 4.325 2.365 ;
        END
        AntennaGateArea 0.2743 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 2.200 2.280 2.360 ;
        RECT  1.990 0.325 2.150 2.360 ;
        RECT  1.375 0.325 1.990 0.485 ;
        RECT  0.760 2.200 1.990 2.360 ;
        RECT  0.295 2.150 0.760 2.360 ;
        END
        AntennaGateArea 0.2847 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 1.455 6.625 1.990 ;
        END
        AntennaGateArea 0.1742 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.515 1.290 1.130 1.580 ;
        END
        AntennaGateArea 0.1885 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 1.280 3.630 1.950 ;
        END
        AntennaGateArea 0.2015 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.700 -0.130 7.380 0.130 ;
        RECT  6.440 -0.130 6.700 0.250 ;
        RECT  4.310 -0.130 6.440 0.130 ;
        RECT  3.370 -0.130 4.310 0.250 ;
        RECT  0.825 -0.130 3.370 0.130 ;
        RECT  0.225 -0.130 0.825 0.340 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 2.740 7.380 3.000 ;
        RECT  6.400 2.170 6.660 3.000 ;
        RECT  3.940 2.740 6.400 3.000 ;
        RECT  3.340 2.570 3.940 3.000 ;
        RECT  0.785 2.740 3.340 3.000 ;
        RECT  0.185 2.570 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.665 0.430 6.865 1.265 ;
        RECT  5.495 0.430 6.665 0.590 ;
        RECT  6.070 0.770 6.145 0.930 ;
        RECT  5.910 0.770 6.070 2.145 ;
        RECT  5.885 0.770 5.910 0.930 ;
        RECT  5.855 1.885 5.910 2.145 ;
        RECT  5.335 0.430 5.495 0.780 ;
        RECT  5.175 0.430 5.335 1.875 ;
        RECT  4.840 1.715 5.175 1.875 ;
        RECT  4.660 0.430 4.880 0.775 ;
        RECT  4.500 0.430 4.660 1.875 ;
        RECT  2.490 0.430 4.500 0.590 ;
        RECT  4.330 1.715 4.500 1.875 ;
        RECT  4.150 0.780 4.320 1.440 ;
        RECT  3.990 0.780 4.150 1.900 ;
        RECT  3.940 0.780 3.990 0.940 ;
        RECT  3.820 1.740 3.990 1.900 ;
        RECT  2.830 0.770 3.080 0.930 ;
        RECT  2.830 1.780 3.020 2.380 ;
        RECT  2.670 0.770 2.830 2.380 ;
        RECT  2.330 0.430 2.490 1.925 ;
        RECT  1.650 0.705 1.810 1.975 ;
        RECT  1.075 1.815 1.650 1.975 ;
        RECT  1.310 0.940 1.470 1.515 ;
        RECT  0.385 0.940 1.310 1.100 ;
        RECT  0.335 0.705 0.385 1.100 ;
        RECT  0.175 0.705 0.335 1.945 ;
        RECT  0.125 0.705 0.175 0.965 ;
        RECT  0.135 1.685 0.175 1.945 ;
    END
END MX3X2MTH

MACRO MX3X4MTH
    CLASS CORE ;
    FOREIGN MX3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.225 0.880 7.280 1.580 ;
        RECT  7.045 0.485 7.225 2.495 ;
        RECT  6.915 0.485 7.045 0.745 ;
        RECT  6.895 1.895 7.045 2.495 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.560 1.115 5.650 1.375 ;
        RECT  5.400 1.115 5.560 2.335 ;
        RECT  4.485 2.175 5.400 2.335 ;
        RECT  3.765 2.150 4.485 2.385 ;
        END
        AntennaGateArea 0.2873 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 2.200 2.280 2.360 ;
        RECT  1.990 0.325 2.150 2.360 ;
        RECT  1.375 0.325 1.990 0.485 ;
        RECT  0.760 2.200 1.990 2.360 ;
        RECT  0.295 2.150 0.760 2.360 ;
        END
        AntennaGateArea 0.2847 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.405 1.700 6.460 1.990 ;
        RECT  6.170 1.345 6.405 1.990 ;
        END
        AntennaGateArea 0.1794 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.525 1.290 1.130 1.580 ;
        END
        AntennaGateArea 0.1885 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.200 1.290 3.590 1.990 ;
        RECT  3.140 1.290 3.200 1.550 ;
        END
        AntennaGateArea 0.2015 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 -0.130 7.790 0.130 ;
        RECT  7.405 -0.130 7.665 0.730 ;
        RECT  6.585 -0.130 7.405 0.130 ;
        RECT  6.325 -0.130 6.585 0.250 ;
        RECT  4.310 -0.130 6.325 0.130 ;
        RECT  3.370 -0.130 4.310 0.250 ;
        RECT  0.825 -0.130 3.370 0.130 ;
        RECT  0.225 -0.130 0.825 0.340 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 2.740 7.790 3.000 ;
        RECT  7.405 1.915 7.665 3.000 ;
        RECT  6.610 2.740 7.405 3.000 ;
        RECT  6.350 2.170 6.610 3.000 ;
        RECT  3.940 2.740 6.350 3.000 ;
        RECT  3.340 2.570 3.940 3.000 ;
        RECT  0.785 2.740 3.340 3.000 ;
        RECT  0.185 2.570 0.785 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.725 0.930 6.865 1.495 ;
        RECT  6.625 0.430 6.725 1.495 ;
        RECT  6.565 0.430 6.625 1.235 ;
        RECT  5.425 0.430 6.565 0.590 ;
        RECT  5.990 0.770 6.075 0.930 ;
        RECT  5.830 0.770 5.990 2.145 ;
        RECT  5.785 0.770 5.830 0.930 ;
        RECT  5.740 1.885 5.830 2.145 ;
        RECT  5.220 0.430 5.425 0.780 ;
        RECT  5.060 0.430 5.220 1.925 ;
        RECT  4.810 1.665 5.060 1.925 ;
        RECT  4.600 0.430 4.880 0.775 ;
        RECT  4.440 0.430 4.600 1.875 ;
        RECT  2.490 0.430 4.440 0.590 ;
        RECT  4.250 1.715 4.440 1.875 ;
        RECT  4.170 1.180 4.260 1.440 ;
        RECT  3.950 0.775 4.170 1.440 ;
        RECT  3.790 0.775 3.950 1.965 ;
        RECT  2.830 0.770 3.080 0.930 ;
        RECT  2.830 1.780 3.020 2.380 ;
        RECT  2.670 0.770 2.830 2.380 ;
        RECT  2.330 0.430 2.490 1.925 ;
        RECT  1.650 0.695 1.810 1.975 ;
        RECT  1.075 1.815 1.650 1.975 ;
        RECT  1.310 0.940 1.470 1.515 ;
        RECT  0.385 0.940 1.310 1.100 ;
        RECT  0.335 0.695 0.385 1.100 ;
        RECT  0.175 0.695 0.335 1.945 ;
        RECT  0.125 0.695 0.175 0.955 ;
        RECT  0.135 1.685 0.175 1.945 ;
    END
END MX3X4MTH

MACRO MX3X8MTH
    CLASS CORE ;
    FOREIGN MX3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.565 0.375 7.675 1.085 ;
        RECT  7.415 0.375 7.565 2.385 ;
        RECT  7.305 0.785 7.415 2.385 ;
        RECT  7.035 0.785 7.305 2.135 ;
        RECT  6.725 0.785 7.035 1.085 ;
        RECT  6.635 1.785 7.035 2.135 ;
        RECT  6.525 0.475 6.725 1.085 ;
        RECT  6.375 1.785 6.635 2.315 ;
        RECT  6.375 0.475 6.525 0.735 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.230 1.005 5.255 1.265 ;
        RECT  5.175 1.005 5.230 1.580 ;
        RECT  5.015 1.005 5.175 2.335 ;
        RECT  3.660 2.175 5.015 2.335 ;
        END
        AntennaGateArea 0.2678 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.675 2.280 2.115 2.440 ;
        RECT  0.675 1.245 0.720 1.580 ;
        RECT  0.515 1.245 0.675 2.440 ;
        RECT  0.430 1.245 0.515 1.580 ;
        END
        AntennaGateArea 0.2821 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.005 1.700 6.050 1.990 ;
        RECT  5.775 1.255 6.005 1.990 ;
        END
        AntennaGateArea 0.182 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 1.230 1.225 1.760 ;
        END
        AntennaGateArea 0.1664 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.110 3.180 1.580 ;
        END
        AntennaGateArea 0.2002 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.165 -0.130 8.200 0.130 ;
        RECT  6.905 -0.130 7.165 0.605 ;
        RECT  3.695 -0.130 6.905 0.130 ;
        RECT  3.095 -0.130 3.695 0.250 ;
        RECT  0.925 -0.130 3.095 0.130 ;
        RECT  0.665 -0.130 0.925 0.710 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 2.740 8.200 3.000 ;
        RECT  7.815 1.800 8.075 3.000 ;
        RECT  6.100 2.740 7.815 3.000 ;
        RECT  5.840 2.185 6.100 3.000 ;
        RECT  3.435 2.740 5.840 3.000 ;
        RECT  3.175 2.520 3.435 3.000 ;
        RECT  0.795 2.740 3.175 3.000 ;
        RECT  0.195 2.620 0.795 3.000 ;
        RECT  0.000 2.740 0.195 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.345 1.305 6.805 1.505 ;
        RECT  6.185 0.915 6.345 1.505 ;
        RECT  5.935 0.915 6.185 1.075 ;
        RECT  5.775 0.310 5.935 1.075 ;
        RECT  4.905 0.310 5.775 0.470 ;
        RECT  5.435 0.665 5.595 2.505 ;
        RECT  5.225 0.665 5.435 0.825 ;
        RECT  5.355 2.245 5.435 2.505 ;
        RECT  4.805 0.310 4.905 0.715 ;
        RECT  4.645 0.310 4.805 1.965 ;
        RECT  4.235 0.390 4.395 1.915 ;
        RECT  4.135 0.390 4.235 0.990 ;
        RECT  4.085 1.755 4.235 1.915 ;
        RECT  2.245 0.430 4.135 0.590 ;
        RECT  3.885 1.195 3.980 1.455 ;
        RECT  3.845 0.770 3.885 1.455 ;
        RECT  3.685 0.770 3.845 1.895 ;
        RECT  3.625 0.770 3.685 1.025 ;
        RECT  3.575 1.735 3.685 1.895 ;
        RECT  2.625 1.790 2.885 2.390 ;
        RECT  2.585 0.770 2.805 0.930 ;
        RECT  2.585 1.790 2.625 1.950 ;
        RECT  2.425 0.770 2.585 1.950 ;
        RECT  2.085 0.385 2.245 2.035 ;
        RECT  1.745 0.525 1.905 2.100 ;
        RECT  1.675 0.525 1.745 0.685 ;
        RECT  1.085 1.940 1.745 2.100 ;
        RECT  1.415 0.425 1.675 0.685 ;
        RECT  1.405 0.890 1.565 1.655 ;
        RECT  0.385 0.890 1.405 1.050 ;
        RECT  0.250 0.765 0.385 1.050 ;
        RECT  0.250 1.800 0.335 2.060 ;
        RECT  0.125 0.765 0.250 2.060 ;
        RECT  0.090 0.890 0.125 2.060 ;
    END
END MX3X8MTH

MACRO MX3XLMTH
    CLASS CORE ;
    FOREIGN MX3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 1.290 6.050 1.580 ;
        RECT  5.825 0.770 6.025 2.025 ;
        RECT  5.765 0.770 5.825 1.005 ;
        RECT  5.765 1.865 5.825 2.025 ;
        END
        AntennaDiffArea 0.224 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 1.075 3.255 1.530 ;
        RECT  2.970 1.075 3.180 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.075 0.515 2.510 ;
        END
        AntennaGateArea 0.1586 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.325 1.290 5.640 1.580 ;
        RECT  5.165 1.145 5.325 1.580 ;
        END
        AntennaGateArea 0.078 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.740 0.920 1.065 1.345 ;
        RECT  0.470 0.920 0.740 1.130 ;
        END
        AntennaGateArea 0.0897 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 1.075 2.790 1.580 ;
        RECT  2.455 1.255 2.570 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.485 -0.130 6.150 0.130 ;
        RECT  4.885 -0.130 5.485 0.250 ;
        RECT  0.925 -0.130 4.885 0.130 ;
        RECT  0.665 -0.130 0.925 0.740 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.945 2.740 6.150 3.000 ;
        RECT  5.345 2.365 5.945 3.000 ;
        RECT  4.720 2.740 5.345 3.000 ;
        RECT  4.120 2.550 4.720 3.000 ;
        RECT  3.445 2.740 4.120 3.000 ;
        RECT  2.845 2.550 3.445 3.000 ;
        RECT  0.955 2.740 2.845 3.000 ;
        RECT  0.695 1.865 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.665 0.375 5.925 0.590 ;
        RECT  4.505 0.430 5.665 0.590 ;
        RECT  4.955 0.770 5.065 0.930 ;
        RECT  4.955 1.935 5.065 2.095 ;
        RECT  4.795 0.770 4.955 2.095 ;
        RECT  4.345 0.430 4.505 2.145 ;
        RECT  3.995 0.770 4.045 0.930 ;
        RECT  3.945 0.770 3.995 2.365 ;
        RECT  3.835 0.395 3.945 2.365 ;
        RECT  3.785 0.395 3.835 0.930 ;
        RECT  1.755 2.205 3.835 2.365 ;
        RECT  2.015 0.395 3.785 0.555 ;
        RECT  3.595 1.075 3.645 1.335 ;
        RECT  3.435 0.735 3.595 2.015 ;
        RECT  3.275 0.735 3.435 0.895 ;
        RECT  3.325 1.755 3.435 2.015 ;
        RECT  2.385 0.735 2.555 0.895 ;
        RECT  2.275 1.760 2.555 1.920 ;
        RECT  2.275 0.735 2.385 1.075 ;
        RECT  2.225 0.735 2.275 1.920 ;
        RECT  2.115 0.915 2.225 1.920 ;
        RECT  1.855 0.395 2.015 0.735 ;
        RECT  1.775 0.975 1.935 2.025 ;
        RECT  1.755 0.575 1.855 0.735 ;
        RECT  1.455 0.975 1.775 1.135 ;
        RECT  1.215 1.865 1.775 2.025 ;
        RECT  1.435 1.315 1.595 1.685 ;
        RECT  1.295 0.525 1.455 1.135 ;
        RECT  0.385 1.525 1.435 1.685 ;
        RECT  0.285 0.580 0.385 0.740 ;
        RECT  0.285 1.525 0.385 1.895 ;
        RECT  0.125 0.580 0.285 1.895 ;
    END
END MX3XLMTH

MACRO MX4X1MTH
    CLASS CORE ;
    FOREIGN MX4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.665 1.700 9.740 1.990 ;
        RECT  9.505 0.740 9.665 1.990 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.780 1.160 8.940 2.560 ;
        RECT  8.660 1.160 8.780 1.580 ;
        RECT  6.965 2.400 8.780 2.560 ;
        END
        AntennaGateArea 0.2301 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 2.400 5.345 2.560 ;
        RECT  4.485 0.310 4.745 0.595 ;
        RECT  3.395 0.435 4.485 0.595 ;
        RECT  3.135 0.310 3.395 0.595 ;
        RECT  2.435 0.435 3.135 0.595 ;
        RECT  2.275 0.310 2.435 0.595 ;
        RECT  1.195 0.310 2.275 0.470 ;
        RECT  1.035 0.310 1.195 2.560 ;
        RECT  0.880 2.150 1.035 2.560 ;
        END
        AntennaGateArea 0.4407 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.330 3.040 1.595 ;
        END
        AntennaGateArea 0.1612 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.120 0.455 1.580 ;
        END
        AntennaGateArea 0.1612 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.645 1.185 4.000 1.725 ;
        END
        AntennaGateArea 0.1612 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.205 0.880 6.490 1.445 ;
        END
        AntennaGateArea 0.1612 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.610 -0.130 9.840 0.130 ;
        RECT  9.010 -0.130 9.610 0.255 ;
        RECT  6.905 -0.130 9.010 0.130 ;
        RECT  6.305 -0.130 6.905 0.280 ;
        RECT  3.935 -0.130 6.305 0.130 ;
        RECT  3.675 -0.130 3.935 0.250 ;
        RECT  0.385 -0.130 3.675 0.130 ;
        RECT  0.125 -0.130 0.385 0.850 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.620 2.740 9.840 3.000 ;
        RECT  9.120 2.555 9.620 3.000 ;
        RECT  6.675 2.740 9.120 3.000 ;
        RECT  6.415 2.570 6.675 3.000 ;
        RECT  0.385 2.740 6.415 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.165 0.435 9.325 1.480 ;
        RECT  8.090 0.435 9.165 0.595 ;
        RECT  8.480 0.795 8.760 0.955 ;
        RECT  8.480 1.820 8.600 2.220 ;
        RECT  8.320 0.795 8.480 2.220 ;
        RECT  6.465 2.060 8.320 2.220 ;
        RECT  7.990 1.720 8.140 1.880 ;
        RECT  7.990 0.435 8.090 0.845 ;
        RECT  7.830 0.435 7.990 1.880 ;
        RECT  7.490 0.460 7.650 1.880 ;
        RECT  7.420 0.460 7.490 0.845 ;
        RECT  7.370 1.720 7.490 1.880 ;
        RECT  5.465 0.460 7.420 0.620 ;
        RECT  7.075 1.140 7.310 1.400 ;
        RECT  7.075 0.800 7.120 0.960 ;
        RECT  7.075 1.720 7.120 1.880 ;
        RECT  6.915 0.800 7.075 1.880 ;
        RECT  6.860 0.800 6.915 0.960 ;
        RECT  6.860 1.720 6.915 1.880 ;
        RECT  6.305 2.060 6.465 2.390 ;
        RECT  5.725 2.230 6.305 2.390 ;
        RECT  6.025 1.625 6.125 2.015 ;
        RECT  5.905 0.800 6.025 2.015 ;
        RECT  5.865 0.800 5.905 1.880 ;
        RECT  5.765 0.800 5.865 0.960 ;
        RECT  5.565 2.060 5.725 2.390 ;
        RECT  5.465 1.720 5.575 1.880 ;
        RECT  1.535 2.060 5.565 2.220 ;
        RECT  5.305 0.460 5.465 1.880 ;
        RECT  4.945 0.775 5.105 1.880 ;
        RECT  4.520 0.775 4.945 0.935 ;
        RECT  4.365 1.720 4.945 1.880 ;
        RECT  4.605 1.145 4.765 1.410 ;
        RECT  4.340 1.145 4.605 1.305 ;
        RECT  4.180 0.800 4.340 1.305 ;
        RECT  3.465 0.800 4.180 0.960 ;
        RECT  3.305 0.800 3.465 1.880 ;
        RECT  2.410 0.940 3.305 1.100 ;
        RECT  3.205 1.720 3.305 1.880 ;
        RECT  2.250 0.940 2.410 1.180 ;
        RECT  2.215 1.020 2.250 1.180 ;
        RECT  2.055 1.020 2.215 1.380 ;
        RECT  1.875 1.720 2.125 1.880 ;
        RECT  1.875 0.680 2.095 0.840 ;
        RECT  1.715 0.680 1.875 1.880 ;
        RECT  1.375 0.750 1.535 2.220 ;
        RECT  0.695 0.750 0.855 1.945 ;
    END
END MX4X1MTH

MACRO MX4X2MTH
    CLASS CORE ;
    FOREIGN MX4X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.125 1.700 10.150 1.990 ;
        RECT  10.075 0.415 10.125 1.015 ;
        RECT  10.075 1.700 10.125 2.400 ;
        RECT  9.915 0.415 10.075 2.400 ;
        RECT  9.865 0.415 9.915 1.015 ;
        RECT  9.865 1.800 9.915 2.400 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.280 1.700 9.335 2.285 ;
        RECT  9.150 1.160 9.280 2.285 ;
        RECT  9.120 1.160 9.150 2.560 ;
        RECT  8.990 1.160 9.120 1.420 ;
        RECT  8.990 2.125 9.120 2.560 ;
        RECT  7.270 2.400 8.990 2.560 ;
        END
        AntennaGateArea 0.2886 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 2.400 5.420 2.560 ;
        RECT  4.745 0.390 5.005 0.595 ;
        RECT  3.965 0.435 4.745 0.595 ;
        RECT  3.705 0.310 3.965 0.595 ;
        RECT  2.725 0.435 3.705 0.595 ;
        RECT  2.565 0.310 2.725 0.595 ;
        RECT  1.195 0.310 2.565 0.470 ;
        RECT  1.035 0.310 1.195 2.560 ;
        RECT  0.880 2.150 1.035 2.360 ;
        END
        AntennaGateArea 0.5759 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.290 3.180 1.580 ;
        RECT  2.705 1.365 2.930 1.580 ;
        RECT  2.585 1.365 2.705 1.525 ;
        END
        AntennaGateArea 0.2028 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.135 0.515 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.185 4.105 1.610 ;
        END
        AntennaGateArea 0.2041 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 0.880 6.870 1.445 ;
        RECT  6.400 1.185 6.565 1.445 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.585 -0.130 10.250 0.130 ;
        RECT  9.325 -0.130 9.585 0.255 ;
        RECT  7.215 -0.130 9.325 0.130 ;
        RECT  6.615 -0.130 7.215 0.255 ;
        RECT  3.165 -0.130 6.615 0.130 ;
        RECT  2.905 -0.130 3.165 0.250 ;
        RECT  0.385 -0.130 2.905 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.585 2.740 10.250 3.000 ;
        RECT  9.325 2.620 9.585 3.000 ;
        RECT  6.955 2.740 9.325 3.000 ;
        RECT  6.695 2.570 6.955 3.000 ;
        RECT  0.385 2.740 6.695 3.000 ;
        RECT  0.125 1.895 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.635 1.220 9.735 1.480 ;
        RECT  9.475 0.435 9.635 1.480 ;
        RECT  8.465 0.435 9.475 0.595 ;
        RECT  8.810 0.795 9.075 0.955 ;
        RECT  8.810 1.670 8.930 1.930 ;
        RECT  8.650 0.795 8.810 2.220 ;
        RECT  6.790 2.060 8.650 2.220 ;
        RECT  8.305 0.435 8.465 1.880 ;
        RECT  8.205 1.720 8.305 1.880 ;
        RECT  7.845 0.395 8.005 1.880 ;
        RECT  5.725 0.435 7.845 0.595 ;
        RECT  7.680 1.720 7.845 1.880 ;
        RECT  7.285 1.160 7.665 1.420 ;
        RECT  7.285 1.720 7.420 1.880 ;
        RECT  7.285 0.800 7.390 0.960 ;
        RECT  7.125 0.800 7.285 1.880 ;
        RECT  6.630 2.060 6.790 2.390 ;
        RECT  5.770 2.230 6.630 2.390 ;
        RECT  6.220 1.805 6.395 1.965 ;
        RECT  6.220 0.795 6.335 0.955 ;
        RECT  6.060 0.795 6.220 1.965 ;
        RECT  5.610 2.060 5.770 2.390 ;
        RECT  5.615 1.720 5.765 1.880 ;
        RECT  5.615 0.435 5.725 0.835 ;
        RECT  5.455 0.435 5.615 1.880 ;
        RECT  1.535 2.060 5.610 2.220 ;
        RECT  5.175 0.775 5.225 0.935 ;
        RECT  5.015 0.775 5.175 1.880 ;
        RECT  4.625 0.775 5.015 0.935 ;
        RECT  4.360 1.720 5.015 1.880 ;
        RECT  4.675 1.150 4.835 1.510 ;
        RECT  4.445 1.150 4.675 1.310 ;
        RECT  4.285 0.800 4.445 1.310 ;
        RECT  3.520 0.800 4.285 0.960 ;
        RECT  3.520 1.720 3.585 1.880 ;
        RECT  3.360 0.800 3.520 1.880 ;
        RECT  2.545 0.800 3.360 0.960 ;
        RECT  3.325 1.720 3.360 1.880 ;
        RECT  2.385 0.800 2.545 1.180 ;
        RECT  1.875 1.720 2.475 1.880 ;
        RECT  2.285 1.020 2.385 1.180 ;
        RECT  2.125 1.020 2.285 1.490 ;
        RECT  1.875 0.680 2.095 0.840 ;
        RECT  1.715 0.680 1.875 1.880 ;
        RECT  1.375 0.750 1.535 2.220 ;
        RECT  0.695 0.400 0.855 1.945 ;
    END
END MX4X2MTH

MACRO MX4X4MTH
    CLASS CORE ;
    FOREIGN MX4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.330 0.785 10.510 1.980 ;
        RECT  10.080 0.785 10.330 0.965 ;
        RECT  10.150 1.800 10.330 1.980 ;
        RECT  9.860 1.800 10.150 2.400 ;
        RECT  9.820 0.365 10.080 0.965 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.280 2.110 9.330 2.400 ;
        RECT  9.150 1.135 9.280 2.400 ;
        RECT  9.120 1.135 9.150 2.560 ;
        RECT  8.990 1.135 9.120 1.395 ;
        RECT  8.990 2.240 9.120 2.560 ;
        RECT  7.290 2.400 8.990 2.560 ;
        END
        AntennaGateArea 0.2886 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 2.400 5.540 2.560 ;
        RECT  4.795 0.390 5.055 0.590 ;
        RECT  2.725 0.430 4.795 0.590 ;
        RECT  2.565 0.310 2.725 0.590 ;
        RECT  1.245 0.310 2.565 0.470 ;
        RECT  1.085 0.310 1.245 2.560 ;
        RECT  0.920 2.110 1.085 2.560 ;
        END
        AntennaGateArea 0.5759 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.290 3.180 1.580 ;
        RECT  2.885 1.365 2.970 1.580 ;
        RECT  2.585 1.365 2.885 1.525 ;
        END
        AntennaGateArea 0.2028 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.180 0.515 1.545 ;
        RECT  0.100 0.880 0.335 1.545 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.185 4.080 1.610 ;
        END
        AntennaGateArea 0.2041 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 0.880 6.870 1.445 ;
        RECT  6.400 1.185 6.565 1.445 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.540 -0.130 10.660 0.130 ;
        RECT  9.280 -0.130 9.540 0.255 ;
        RECT  7.215 -0.130 9.280 0.130 ;
        RECT  6.615 -0.130 7.215 0.255 ;
        RECT  3.215 -0.130 6.615 0.130 ;
        RECT  2.955 -0.130 3.215 0.250 ;
        RECT  0.390 -0.130 2.955 0.130 ;
        RECT  0.130 -0.130 0.390 0.605 ;
        RECT  0.125 -0.130 0.130 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.580 2.740 10.660 3.000 ;
        RECT  9.320 2.620 9.580 3.000 ;
        RECT  6.955 2.740 9.320 3.000 ;
        RECT  6.695 2.570 6.955 3.000 ;
        RECT  0.390 2.740 6.695 3.000 ;
        RECT  0.130 1.815 0.390 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.625 1.215 10.150 1.475 ;
        RECT  9.465 0.435 9.625 1.475 ;
        RECT  8.470 0.435 9.465 0.595 ;
        RECT  8.810 0.795 9.090 0.955 ;
        RECT  8.810 1.795 8.930 2.055 ;
        RECT  8.650 0.795 8.810 2.220 ;
        RECT  6.790 2.060 8.650 2.220 ;
        RECT  8.310 0.435 8.470 1.880 ;
        RECT  8.210 1.720 8.310 1.880 ;
        RECT  8.000 0.395 8.070 0.995 ;
        RECT  7.840 0.395 8.000 1.880 ;
        RECT  7.810 0.395 7.840 0.995 ;
        RECT  7.670 1.720 7.840 1.880 ;
        RECT  5.825 0.435 7.810 0.595 ;
        RECT  7.320 1.175 7.660 1.435 ;
        RECT  7.320 0.775 7.560 0.935 ;
        RECT  7.320 1.720 7.420 1.880 ;
        RECT  7.160 0.775 7.320 1.880 ;
        RECT  6.630 2.060 6.790 2.390 ;
        RECT  5.880 2.230 6.630 2.390 ;
        RECT  6.220 1.805 6.445 1.965 ;
        RECT  6.220 0.795 6.335 0.955 ;
        RECT  6.060 0.795 6.220 1.965 ;
        RECT  5.720 2.060 5.880 2.390 ;
        RECT  5.720 0.435 5.825 0.840 ;
        RECT  5.560 0.435 5.720 1.880 ;
        RECT  1.585 2.060 5.720 2.220 ;
        RECT  5.460 1.720 5.560 1.880 ;
        RECT  5.225 0.775 5.275 0.935 ;
        RECT  5.065 0.775 5.225 1.880 ;
        RECT  4.675 0.775 5.065 0.935 ;
        RECT  4.480 1.720 5.065 1.880 ;
        RECT  4.725 1.150 4.885 1.465 ;
        RECT  4.420 1.150 4.725 1.310 ;
        RECT  4.260 0.800 4.420 1.310 ;
        RECT  3.580 0.800 4.260 0.960 ;
        RECT  3.580 1.720 3.615 1.880 ;
        RECT  3.420 0.800 3.580 1.880 ;
        RECT  2.690 0.950 3.420 1.110 ;
        RECT  3.355 1.720 3.420 1.880 ;
        RECT  2.530 0.950 2.690 1.180 ;
        RECT  2.285 1.020 2.530 1.180 ;
        RECT  1.925 1.720 2.475 1.880 ;
        RECT  1.925 0.680 2.355 0.840 ;
        RECT  2.125 1.020 2.285 1.425 ;
        RECT  1.765 0.680 1.925 1.880 ;
        RECT  1.425 0.750 1.585 2.220 ;
        RECT  0.855 0.400 0.905 1.000 ;
        RECT  0.855 1.735 0.905 1.895 ;
        RECT  0.695 0.400 0.855 1.895 ;
        RECT  0.645 0.400 0.695 1.000 ;
        RECT  0.645 1.735 0.695 1.895 ;
    END
END MX4X4MTH

MACRO MX4X8MTH
    CLASS CORE ;
    FOREIGN MX4X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.930 0.410 11.300 2.400 ;
        RECT  10.305 1.290 10.930 1.640 ;
        RECT  9.975 0.405 10.305 2.405 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.280 1.700 9.330 1.990 ;
        RECT  9.160 1.160 9.280 2.405 ;
        RECT  9.120 1.160 9.160 2.560 ;
        RECT  9.000 1.160 9.120 1.420 ;
        RECT  9.000 2.245 9.120 2.560 ;
        RECT  7.340 2.400 9.000 2.560 ;
        END
        AntennaGateArea 0.2886 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.245 2.400 5.605 2.560 ;
        RECT  4.795 0.390 5.055 0.590 ;
        RECT  2.660 0.430 4.795 0.590 ;
        RECT  2.500 0.310 2.660 0.590 ;
        RECT  1.245 0.310 2.500 0.470 ;
        RECT  1.085 0.310 1.245 2.560 ;
        RECT  0.920 2.110 1.085 2.560 ;
        END
        AntennaGateArea 0.5759 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.290 3.180 1.580 ;
        RECT  2.655 1.365 2.970 1.580 ;
        RECT  2.585 1.365 2.655 1.525 ;
        END
        AntennaGateArea 0.2028 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.120 0.515 1.485 ;
        RECT  0.100 0.880 0.335 1.485 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.185 4.195 1.610 ;
        END
        AntennaGateArea 0.2041 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.565 0.880 6.870 1.445 ;
        RECT  6.465 1.185 6.565 1.445 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 -0.130 11.890 0.130 ;
        RECT  11.505 -0.130 11.765 0.960 ;
        RECT  10.745 -0.130 11.505 0.130 ;
        RECT  10.485 -0.130 10.745 0.960 ;
        RECT  9.695 -0.130 10.485 0.130 ;
        RECT  9.435 -0.130 9.695 0.250 ;
        RECT  7.555 -0.130 9.435 0.130 ;
        RECT  6.615 -0.130 7.555 0.250 ;
        RECT  3.215 -0.130 6.615 0.130 ;
        RECT  2.955 -0.130 3.215 0.250 ;
        RECT  0.385 -0.130 2.955 0.130 ;
        RECT  0.125 -0.130 0.385 0.605 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 2.740 11.890 3.000 ;
        RECT  11.505 1.800 11.765 3.000 ;
        RECT  10.745 2.740 11.505 3.000 ;
        RECT  10.485 1.915 10.745 3.000 ;
        RECT  9.715 2.740 10.485 3.000 ;
        RECT  9.515 1.800 9.715 3.000 ;
        RECT  9.435 2.570 9.515 3.000 ;
        RECT  6.990 2.740 9.435 3.000 ;
        RECT  6.730 2.570 6.990 3.000 ;
        RECT  0.385 2.740 6.730 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.595 0.435 9.755 1.480 ;
        RECT  8.455 0.435 9.595 0.595 ;
        RECT  8.820 0.795 9.185 0.955 ;
        RECT  8.820 1.795 8.940 2.055 ;
        RECT  8.660 0.795 8.820 2.220 ;
        RECT  6.790 2.060 8.660 2.220 ;
        RECT  8.455 1.720 8.480 1.880 ;
        RECT  8.295 0.435 8.455 1.880 ;
        RECT  8.220 1.720 8.295 1.880 ;
        RECT  8.040 0.395 8.115 0.995 ;
        RECT  7.955 0.395 8.040 1.880 ;
        RECT  7.880 0.435 7.955 1.880 ;
        RECT  5.825 0.435 7.880 0.595 ;
        RECT  7.710 1.720 7.880 1.880 ;
        RECT  7.300 1.180 7.700 1.440 ;
        RECT  7.300 0.775 7.610 0.935 ;
        RECT  7.300 1.720 7.460 1.880 ;
        RECT  7.140 0.775 7.300 1.880 ;
        RECT  6.630 2.060 6.790 2.390 ;
        RECT  5.945 2.230 6.630 2.390 ;
        RECT  6.285 1.805 6.450 1.965 ;
        RECT  6.285 0.795 6.335 0.955 ;
        RECT  6.125 0.795 6.285 1.965 ;
        RECT  6.075 0.795 6.125 0.955 ;
        RECT  5.785 2.060 5.945 2.390 ;
        RECT  5.720 0.435 5.825 0.840 ;
        RECT  1.585 2.060 5.785 2.220 ;
        RECT  5.560 0.435 5.720 1.880 ;
        RECT  5.460 1.720 5.560 1.880 ;
        RECT  5.280 0.775 5.315 0.935 ;
        RECT  5.120 0.775 5.280 1.880 ;
        RECT  4.715 0.775 5.120 0.935 ;
        RECT  4.545 1.720 5.120 1.880 ;
        RECT  4.780 1.150 4.940 1.410 ;
        RECT  4.535 1.150 4.780 1.310 ;
        RECT  4.375 0.800 4.535 1.310 ;
        RECT  3.610 0.800 4.375 0.960 ;
        RECT  3.610 1.720 3.640 1.880 ;
        RECT  3.450 0.800 3.610 1.880 ;
        RECT  2.645 0.935 3.450 1.095 ;
        RECT  3.330 1.720 3.450 1.880 ;
        RECT  2.485 0.935 2.645 1.180 ;
        RECT  2.285 1.020 2.485 1.180 ;
        RECT  1.925 1.720 2.475 1.880 ;
        RECT  2.125 1.020 2.285 1.425 ;
        RECT  1.925 0.680 2.215 0.840 ;
        RECT  1.765 0.680 1.925 1.880 ;
        RECT  1.425 0.750 1.585 2.220 ;
        RECT  0.855 1.735 0.905 1.895 ;
        RECT  0.695 0.400 0.855 1.895 ;
        RECT  0.645 1.735 0.695 1.895 ;
    END
END MX4X8MTH

MACRO MX4XLMTH
    CLASS CORE ;
    FOREIGN MX4XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.665 1.700 9.740 1.990 ;
        RECT  9.505 0.740 9.665 1.990 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.775 1.160 8.935 2.560 ;
        RECT  8.710 1.160 8.775 1.580 ;
        RECT  7.495 2.400 8.775 2.560 ;
        RECT  8.625 1.160 8.710 1.420 ;
        END
        AntennaGateArea 0.143 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.195 2.400 5.775 2.560 ;
        RECT  4.805 0.370 5.065 0.595 ;
        RECT  3.355 0.435 4.805 0.595 ;
        RECT  3.095 0.340 3.355 0.595 ;
        RECT  2.465 0.435 3.095 0.595 ;
        RECT  2.305 0.310 2.465 0.595 ;
        RECT  1.195 0.310 2.305 0.470 ;
        RECT  1.035 0.310 1.195 2.560 ;
        RECT  0.880 2.150 1.035 2.360 ;
        END
        AntennaGateArea 0.2548 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 1.330 3.220 1.540 ;
        RECT  2.560 1.330 3.040 1.595 ;
        RECT  2.485 1.435 2.560 1.595 ;
        END
        AntennaGateArea 0.0897 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.210 0.515 1.580 ;
        END
        AntennaGateArea 0.0897 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.740 1.185 4.055 1.700 ;
        END
        AntennaGateArea 0.0897 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.250 0.880 6.460 1.445 ;
        RECT  6.185 1.185 6.250 1.445 ;
        END
        AntennaGateArea 0.0897 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.575 -0.130 9.840 0.130 ;
        RECT  8.975 -0.130 9.575 0.255 ;
        RECT  8.485 -0.130 8.975 0.130 ;
        RECT  7.885 -0.130 8.485 0.255 ;
        RECT  4.405 -0.130 7.885 0.130 ;
        RECT  3.805 -0.130 4.405 0.250 ;
        RECT  2.915 -0.130 3.805 0.130 ;
        RECT  2.655 -0.130 2.915 0.250 ;
        RECT  0.725 -0.130 2.655 0.130 ;
        RECT  0.385 -0.130 0.725 0.450 ;
        RECT  0.125 -0.130 0.385 1.010 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.615 2.740 9.840 3.000 ;
        RECT  9.115 2.295 9.615 3.000 ;
        RECT  6.995 2.740 9.115 3.000 ;
        RECT  6.395 2.415 6.995 3.000 ;
        RECT  0.725 2.740 6.395 3.000 ;
        RECT  0.385 2.540 0.725 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.165 0.435 9.325 1.480 ;
        RECT  8.105 0.435 9.165 0.595 ;
        RECT  8.445 0.795 8.725 0.955 ;
        RECT  8.445 1.750 8.595 2.220 ;
        RECT  8.285 0.795 8.445 2.220 ;
        RECT  1.535 2.060 8.285 2.220 ;
        RECT  7.945 0.435 8.105 1.880 ;
        RECT  7.815 1.720 7.945 1.880 ;
        RECT  7.470 0.330 7.630 1.880 ;
        RECT  7.405 0.330 7.470 0.845 ;
        RECT  7.335 1.720 7.470 1.880 ;
        RECT  5.445 0.330 7.405 0.490 ;
        RECT  7.105 0.990 7.240 1.250 ;
        RECT  7.085 0.670 7.105 1.250 ;
        RECT  6.925 0.670 7.085 1.880 ;
        RECT  6.845 0.670 6.925 0.830 ;
        RECT  6.825 1.720 6.925 1.880 ;
        RECT  6.005 1.720 6.115 1.880 ;
        RECT  5.845 0.795 6.005 1.880 ;
        RECT  5.745 0.795 5.845 0.955 ;
        RECT  5.445 1.720 5.575 1.880 ;
        RECT  5.285 0.330 5.445 1.880 ;
        RECT  5.225 0.750 5.285 1.010 ;
        RECT  4.885 0.800 5.045 1.880 ;
        RECT  4.605 0.800 4.885 0.960 ;
        RECT  4.405 1.720 4.885 1.880 ;
        RECT  4.545 1.145 4.705 1.410 ;
        RECT  4.425 1.145 4.545 1.305 ;
        RECT  4.265 0.800 4.425 1.305 ;
        RECT  3.560 0.800 4.265 0.960 ;
        RECT  3.400 0.800 3.560 1.880 ;
        RECT  3.295 0.800 3.400 1.100 ;
        RECT  3.205 1.720 3.400 1.880 ;
        RECT  2.385 0.940 3.295 1.100 ;
        RECT  2.225 0.940 2.385 1.250 ;
        RECT  2.215 1.090 2.225 1.250 ;
        RECT  2.055 1.090 2.215 1.380 ;
        RECT  1.875 1.720 2.125 1.880 ;
        RECT  1.875 0.650 2.045 0.910 ;
        RECT  1.715 0.650 1.875 1.880 ;
        RECT  1.375 0.650 1.535 2.220 ;
        RECT  0.695 0.750 0.855 1.970 ;
    END
END MX4XLMTH

MACRO MXI2DX1MTH
    CLASS CORE ;
    FOREIGN MXI2DX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.840 0.710 4.000 2.005 ;
        RECT  3.715 0.710 3.840 0.970 ;
        RECT  3.715 1.700 3.840 2.005 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.535 1.580 ;
        END
        AntennaGateArea 0.0689 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.835 0.520 1.995 2.005 ;
        RECT  1.785 0.520 1.835 0.780 ;
        RECT  1.740 1.700 1.835 2.005 ;
        RECT  1.675 1.745 1.740 2.005 ;
        END
        AntennaDiffArea 0.282 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 0.520 3.015 0.780 ;
        RECT  2.845 1.735 2.955 1.895 ;
        RECT  2.685 0.520 2.845 1.895 ;
        RECT  2.560 1.290 2.685 1.580 ;
        END
        AntennaDiffArea 0.282 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 -0.130 4.100 0.130 ;
        RECT  3.265 -0.130 3.865 0.415 ;
        RECT  0.915 -0.130 3.265 0.130 ;
        RECT  0.315 -0.130 0.915 0.515 ;
        RECT  0.000 -0.130 0.315 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  2.835 2.415 3.435 3.000 ;
        RECT  0.855 2.740 2.835 3.000 ;
        RECT  0.255 2.250 0.855 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.435 1.200 3.610 1.460 ;
        RECT  3.275 1.200 3.435 2.235 ;
        RECT  2.445 2.075 3.275 2.235 ;
        RECT  2.380 0.520 2.505 0.780 ;
        RECT  2.380 1.805 2.445 2.235 ;
        RECT  2.285 0.520 2.380 2.235 ;
        RECT  2.220 0.520 2.285 1.965 ;
        RECT  2.185 1.805 2.220 1.965 ;
        RECT  1.485 2.295 1.775 2.455 ;
        RECT  1.485 0.370 1.595 0.530 ;
        RECT  1.325 0.370 1.485 2.455 ;
        RECT  1.225 0.765 1.325 1.025 ;
        RECT  1.165 1.710 1.325 1.970 ;
        RECT  0.925 1.195 1.085 1.455 ;
        RECT  0.765 0.865 0.925 1.920 ;
        RECT  0.385 0.865 0.765 1.025 ;
        RECT  0.125 1.760 0.765 1.920 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END MXI2DX1MTH

MACRO MXI2DX2MTH
    CLASS CORE ;
    FOREIGN MXI2DX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.925 1.700 4.000 2.410 ;
        RECT  3.925 0.395 3.975 0.995 ;
        RECT  3.765 0.395 3.925 2.410 ;
        RECT  3.715 0.395 3.765 0.995 ;
        RECT  3.715 1.810 3.765 2.410 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.145 0.535 1.580 ;
        END
        AntennaGateArea 0.1066 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.965 1.600 2.005 2.200 ;
        RECT  1.805 0.675 1.965 2.200 ;
        RECT  1.635 0.675 1.805 0.935 ;
        RECT  1.715 1.600 1.805 2.200 ;
        END
        AntennaDiffArea 0.431 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.855 1.745 3.025 1.905 ;
        RECT  2.855 0.490 2.915 0.750 ;
        RECT  2.695 0.490 2.855 1.905 ;
        RECT  2.655 0.490 2.695 1.170 ;
        RECT  2.560 0.880 2.655 1.170 ;
        END
        AntennaDiffArea 0.423 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 -0.130 4.100 0.130 ;
        RECT  3.205 -0.130 3.465 0.970 ;
        RECT  0.815 -0.130 3.205 0.130 ;
        RECT  0.215 -0.130 0.815 0.315 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 2.740 4.100 3.000 ;
        RECT  3.175 2.425 3.435 3.000 ;
        RECT  0.955 2.740 3.175 3.000 ;
        RECT  0.355 2.385 0.955 3.000 ;
        RECT  0.000 2.740 0.355 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.435 1.200 3.580 1.460 ;
        RECT  3.275 1.200 3.435 2.245 ;
        RECT  2.515 2.085 3.275 2.245 ;
        RECT  2.380 1.850 2.515 2.245 ;
        RECT  2.380 0.490 2.405 0.750 ;
        RECT  2.220 0.490 2.380 2.245 ;
        RECT  2.145 0.490 2.220 0.750 ;
        RECT  1.445 2.400 1.865 2.560 ;
        RECT  1.445 0.310 1.525 0.470 ;
        RECT  1.285 0.310 1.445 2.560 ;
        RECT  1.125 0.310 1.285 0.935 ;
        RECT  0.945 1.305 1.040 1.565 ;
        RECT  0.785 0.745 0.945 1.920 ;
        RECT  0.385 0.745 0.785 0.905 ;
        RECT  0.385 1.760 0.785 1.920 ;
        RECT  0.125 0.645 0.385 0.905 ;
        RECT  0.125 1.760 0.385 2.020 ;
    END
END MXI2DX2MTH

MACRO MXI2DX4MTH
    CLASS CORE ;
    FOREIGN MXI2DX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.105 1.270 5.230 1.585 ;
        RECT  4.945 0.395 5.105 2.410 ;
        RECT  4.845 0.395 4.945 0.995 ;
        RECT  4.845 1.810 4.945 2.410 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.535 1.615 ;
        END
        AntennaGateArea 0.2054 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 1.290 2.770 1.620 ;
        RECT  2.450 1.290 2.555 1.880 ;
        RECT  2.290 0.675 2.450 1.880 ;
        RECT  2.185 0.675 2.290 0.935 ;
        END
        AntennaDiffArea 0.506 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.475 0.880 3.590 1.945 ;
        RECT  3.315 0.675 3.475 1.945 ;
        RECT  3.205 0.675 3.315 0.935 ;
        END
        AntennaDiffArea 0.518 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 0.995 ;
        RECT  4.540 -0.130 5.355 0.130 ;
        RECT  4.280 -0.130 4.540 0.980 ;
        RECT  0.000 -0.130 4.280 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 1.800 5.615 3.000 ;
        RECT  4.595 2.740 5.355 3.000 ;
        RECT  4.335 1.800 4.595 3.000 ;
        RECT  0.955 2.740 4.335 3.000 ;
        RECT  0.695 2.230 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.085 1.205 4.760 1.465 ;
        RECT  3.825 1.205 4.085 2.285 ;
        RECT  3.715 0.335 3.975 0.720 ;
        RECT  3.065 2.125 3.825 2.285 ;
        RECT  2.955 0.335 3.715 0.495 ;
        RECT  2.805 1.810 3.065 2.285 ;
        RECT  2.695 0.335 2.955 0.735 ;
        RECT  2.005 2.060 2.805 2.220 ;
        RECT  2.005 0.335 2.695 0.495 ;
        RECT  1.845 0.335 2.005 2.220 ;
        RECT  1.495 2.400 1.870 2.560 ;
        RECT  1.675 0.675 1.845 0.935 ;
        RECT  1.800 1.820 1.845 2.220 ;
        RECT  1.495 0.310 1.665 0.470 ;
        RECT  1.335 0.310 1.495 2.560 ;
        RECT  1.145 0.675 1.335 0.935 ;
        RECT  1.290 1.855 1.335 2.560 ;
        RECT  0.965 1.230 1.110 1.490 ;
        RECT  0.805 0.815 0.965 2.050 ;
        RECT  0.385 0.815 0.805 0.975 ;
        RECT  0.385 1.890 0.805 2.050 ;
        RECT  0.125 0.375 0.385 0.975 ;
        RECT  0.125 1.890 0.385 2.490 ;
    END
END MXI2DX4MTH

MACRO MXI2DX8MTH
    CLASS CORE ;
    FOREIGN MXI2DX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.875 1.210 8.920 2.455 ;
        RECT  8.525 0.425 8.875 2.455 ;
        RECT  7.895 1.210 8.525 1.560 ;
        RECT  7.545 0.395 7.895 2.410 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.405 1.235 0.905 1.615 ;
        END
        AntennaGateArea 0.4108 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.310 1.595 4.410 1.855 ;
        RECT  4.150 0.675 4.310 1.855 ;
        RECT  4.035 0.675 4.150 0.935 ;
        RECT  3.390 1.585 4.150 1.745 ;
        RECT  3.275 1.585 3.390 1.880 ;
        RECT  3.115 0.675 3.275 1.880 ;
        RECT  3.015 0.675 3.115 0.935 ;
        RECT  2.970 1.290 3.115 1.620 ;
        END
        AntennaDiffArea 0.988 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.355 1.765 6.455 2.025 ;
        RECT  6.195 0.675 6.355 2.025 ;
        RECT  6.080 0.675 6.195 1.090 ;
        RECT  5.330 0.930 6.080 1.090 ;
        RECT  5.330 1.770 5.435 2.030 ;
        RECT  5.170 0.675 5.330 2.030 ;
        RECT  5.020 0.675 5.170 1.170 ;
        END
        AntennaDiffArea 1.043 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.255 -0.130 9.430 0.130 ;
        RECT  9.095 -0.130 9.255 0.955 ;
        RECT  8.235 -0.130 9.095 0.130 ;
        RECT  8.075 -0.130 8.235 0.955 ;
        RECT  7.235 -0.130 8.075 0.130 ;
        RECT  6.975 -0.130 7.235 0.300 ;
        RECT  1.325 -0.130 6.975 0.130 ;
        RECT  1.065 -0.130 1.325 0.300 ;
        RECT  0.000 -0.130 1.065 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.335 2.740 9.430 3.000 ;
        RECT  8.175 1.810 8.335 3.000 ;
        RECT  7.335 2.740 8.175 3.000 ;
        RECT  7.075 2.560 7.335 3.000 ;
        RECT  2.025 2.740 7.075 3.000 ;
        RECT  1.085 2.565 2.025 3.000 ;
        RECT  0.000 2.740 1.085 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.965 1.205 7.365 1.465 ;
        RECT  6.705 1.205 6.965 2.370 ;
        RECT  6.750 0.640 6.850 0.900 ;
        RECT  6.590 0.335 6.750 0.900 ;
        RECT  5.945 2.210 6.705 2.370 ;
        RECT  5.830 0.335 6.590 0.495 ;
        RECT  5.685 1.770 5.945 2.370 ;
        RECT  5.570 0.335 5.830 0.750 ;
        RECT  4.920 2.210 5.685 2.370 ;
        RECT  4.805 0.335 5.570 0.495 ;
        RECT  4.660 1.940 4.920 2.370 ;
        RECT  4.545 0.335 4.805 0.735 ;
        RECT  4.655 2.060 4.660 2.370 ;
        RECT  3.900 2.060 4.655 2.220 ;
        RECT  3.785 0.335 4.545 0.495 ;
        RECT  3.640 1.955 3.900 2.220 ;
        RECT  3.525 0.335 3.785 0.750 ;
        RECT  2.845 2.060 3.640 2.220 ;
        RECT  2.835 0.335 3.525 0.495 ;
        RECT  2.785 1.830 2.845 2.220 ;
        RECT  2.785 0.335 2.835 0.935 ;
        RECT  2.675 0.335 2.785 2.220 ;
        RECT  2.375 2.400 2.705 2.560 ;
        RECT  2.625 0.675 2.675 2.220 ;
        RECT  2.555 0.675 2.625 0.935 ;
        RECT  2.585 1.830 2.625 2.220 ;
        RECT  2.375 0.310 2.495 0.470 ;
        RECT  2.215 0.310 2.375 2.560 ;
        RECT  1.725 0.750 2.215 0.910 ;
        RECT  1.810 1.950 2.215 2.110 ;
        RECT  1.280 1.230 1.845 1.490 ;
        RECT  1.550 1.850 1.810 2.110 ;
        RECT  1.465 0.650 1.725 0.910 ;
        RECT  1.120 0.865 1.280 2.065 ;
        RECT  0.785 0.865 1.120 1.025 ;
        RECT  0.785 1.905 1.120 2.065 ;
        RECT  0.525 0.425 0.785 1.025 ;
        RECT  0.525 1.905 0.785 2.505 ;
    END
END MXI2DX8MTH

MACRO MXI2DXLMTH
    CLASS CORE ;
    FOREIGN MXI2DXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.840 0.765 4.000 2.005 ;
        RECT  3.715 0.765 3.840 1.025 ;
        RECT  3.715 1.700 3.840 2.005 ;
        END
        AntennaDiffArea 0.224 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.535 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 0.520 1.985 2.005 ;
        RECT  1.785 0.520 1.825 0.780 ;
        RECT  1.675 1.700 1.825 2.005 ;
        END
        AntennaDiffArea 0.204 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 0.520 3.015 0.780 ;
        RECT  2.845 1.760 2.955 1.920 ;
        RECT  2.685 0.520 2.845 1.920 ;
        RECT  2.560 1.290 2.685 1.580 ;
        END
        AntennaDiffArea 0.204 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 -0.130 4.100 0.130 ;
        RECT  3.265 -0.130 3.865 0.415 ;
        RECT  0.915 -0.130 3.265 0.130 ;
        RECT  0.315 -0.130 0.915 0.515 ;
        RECT  0.000 -0.130 0.315 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 2.740 4.100 3.000 ;
        RECT  3.175 2.440 3.805 3.000 ;
        RECT  0.855 2.740 3.175 3.000 ;
        RECT  0.255 2.220 0.855 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.435 1.205 3.635 1.465 ;
        RECT  3.275 1.205 3.435 2.260 ;
        RECT  2.445 2.100 3.275 2.260 ;
        RECT  2.345 0.520 2.505 0.780 ;
        RECT  2.345 1.760 2.445 2.260 ;
        RECT  2.185 0.520 2.345 2.260 ;
        RECT  1.485 2.295 1.795 2.455 ;
        RECT  1.485 0.370 1.595 0.530 ;
        RECT  1.325 0.370 1.485 2.455 ;
        RECT  1.225 0.765 1.325 1.025 ;
        RECT  1.165 1.710 1.325 1.970 ;
        RECT  0.925 1.205 1.035 1.465 ;
        RECT  0.765 0.865 0.925 1.920 ;
        RECT  0.385 0.865 0.765 1.025 ;
        RECT  0.125 1.760 0.765 1.920 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END MXI2DXLMTH

MACRO MXI2X12MTH
    CLASS CORE ;
    FOREIGN MXI2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.410 1.125 12.855 1.745 ;
        RECT  11.870 0.785 12.410 2.085 ;
        RECT  8.490 0.785 11.870 1.075 ;
        RECT  8.900 1.675 11.870 2.085 ;
        RECT  8.455 1.675 8.900 2.520 ;
        RECT  8.230 0.425 8.490 1.075 ;
        RECT  5.510 2.120 8.455 2.520 ;
        RECT  5.450 0.785 8.230 1.075 ;
        RECT  5.180 0.720 5.450 1.075 ;
        END
        AntennaDiffArea 4.146 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.595 1.290 4.540 1.580 ;
        END
        AntennaGateArea 1.7602 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.585 1.230 15.175 1.580 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 1.235 2.445 1.580 ;
        END
        AntennaGateArea 1.2324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.450 -0.130 15.580 0.130 ;
        RECT  15.190 -0.130 15.450 0.905 ;
        RECT  14.415 -0.130 15.190 0.130 ;
        RECT  14.155 -0.130 14.415 0.565 ;
        RECT  13.375 -0.130 14.155 0.130 ;
        RECT  13.115 -0.130 13.375 0.565 ;
        RECT  2.430 -0.130 13.115 0.130 ;
        RECT  2.170 -0.130 2.430 0.615 ;
        RECT  1.410 -0.130 2.170 0.130 ;
        RECT  1.150 -0.130 1.410 0.615 ;
        RECT  0.390 -0.130 1.150 0.130 ;
        RECT  0.130 -0.130 0.390 0.955 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.450 2.740 15.580 3.000 ;
        RECT  15.190 1.915 15.450 3.000 ;
        RECT  14.415 2.740 15.190 3.000 ;
        RECT  14.155 2.305 14.415 3.000 ;
        RECT  13.375 2.740 14.155 3.000 ;
        RECT  13.115 2.305 13.375 3.000 ;
        RECT  4.450 2.740 13.115 3.000 ;
        RECT  4.190 2.600 4.450 3.000 ;
        RECT  2.425 2.740 4.190 3.000 ;
        RECT  2.165 2.250 2.425 3.000 ;
        RECT  1.405 2.740 2.165 3.000 ;
        RECT  1.145 2.250 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.820 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.675 0.405 14.935 0.905 ;
        RECT  14.675 1.915 14.935 2.515 ;
        RECT  13.895 0.745 14.675 0.905 ;
        RECT  13.895 1.965 14.675 2.125 ;
        RECT  13.635 0.405 13.895 0.905 ;
        RECT  13.635 1.915 13.895 2.515 ;
        RECT  13.405 0.745 13.635 0.905 ;
        RECT  13.405 1.965 13.635 2.125 ;
        RECT  13.245 0.745 13.405 2.125 ;
        RECT  12.855 0.745 13.245 0.905 ;
        RECT  12.855 1.965 13.245 2.125 ;
        RECT  12.595 0.405 12.855 0.905 ;
        RECT  12.595 1.965 12.855 2.465 ;
        RECT  8.740 0.405 12.595 0.565 ;
        RECT  9.080 2.305 12.595 2.465 ;
        RECT  4.990 1.295 11.690 1.455 ;
        RECT  5.330 1.735 8.275 1.895 ;
        RECT  7.680 0.315 7.940 0.565 ;
        RECT  6.920 0.315 7.680 0.475 ;
        RECT  6.660 0.315 6.920 0.565 ;
        RECT  5.900 0.315 6.660 0.475 ;
        RECT  5.640 0.315 5.900 0.565 ;
        RECT  2.940 0.315 5.640 0.475 ;
        RECT  5.170 1.735 5.330 2.335 ;
        RECT  2.940 2.175 5.170 2.335 ;
        RECT  4.810 0.655 4.990 1.930 ;
        RECT  3.680 0.655 4.810 0.815 ;
        RECT  3.650 1.770 4.810 1.930 ;
        RECT  2.780 0.315 2.940 2.420 ;
        RECT  2.680 0.315 2.780 0.955 ;
        RECT  2.675 1.820 2.780 2.420 ;
        RECT  1.920 0.795 2.680 0.955 ;
        RECT  1.915 1.820 2.675 1.980 ;
        RECT  1.660 0.355 1.920 0.955 ;
        RECT  1.655 1.820 1.915 2.420 ;
        RECT  0.900 0.795 1.660 0.955 ;
        RECT  0.895 1.820 1.655 1.980 ;
        RECT  0.640 0.355 0.900 0.955 ;
        RECT  0.635 1.820 0.895 2.420 ;
    END
END MXI2X12MTH

MACRO MXI2X1MTH
    CLASS CORE ;
    FOREIGN MXI2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 2.150 2.400 2.360 ;
        RECT  2.125 1.010 2.265 2.360 ;
        RECT  2.105 0.630 2.125 2.360 ;
        RECT  1.965 0.630 2.105 1.170 ;
        END
        AntennaDiffArea 0.518 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 0.310 1.835 0.470 ;
        RECT  1.575 0.310 1.735 0.635 ;
        RECT  0.720 0.475 1.575 0.635 ;
        RECT  0.560 0.475 0.720 1.580 ;
        RECT  0.430 1.245 0.560 1.580 ;
        END
        AntennaGateArea 0.182 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.155 1.225 1.615 ;
        END
        AntennaGateArea 0.1209 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.290 3.590 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.950 ;
        RECT  2.665 -0.130 3.305 0.285 ;
        RECT  1.085 -0.130 2.665 0.130 ;
        RECT  0.485 -0.130 1.085 0.285 ;
        RECT  0.000 -0.130 0.485 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.365 2.740 3.690 3.000 ;
        RECT  3.105 1.760 3.365 3.000 ;
        RECT  0.905 2.740 3.105 3.000 ;
        RECT  0.745 2.135 0.905 3.000 ;
        RECT  0.000 2.740 0.745 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.775 0.680 3.025 0.840 ;
        RECT  2.615 0.680 2.775 2.100 ;
        RECT  2.425 0.680 2.615 0.840 ;
        RECT  1.765 1.350 1.925 2.415 ;
        RECT  1.245 2.255 1.765 2.415 ;
        RECT  1.585 0.815 1.635 0.975 ;
        RECT  1.425 0.815 1.585 2.075 ;
        RECT  1.375 0.815 1.425 0.975 ;
        RECT  1.085 1.795 1.245 2.415 ;
        RECT  0.385 1.795 1.085 1.955 ;
        RECT  0.250 1.760 0.385 1.955 ;
        RECT  0.250 0.765 0.335 1.025 ;
        RECT  0.090 0.765 0.250 1.955 ;
    END
END MXI2X1MTH

MACRO MXI2X2MTH
    CLASS CORE ;
    FOREIGN MXI2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.590 2.925 2.400 ;
        RECT  2.365 1.590 2.560 1.750 ;
        RECT  2.205 0.765 2.365 1.750 ;
        END
        AntennaDiffArea 0.654 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 1.150 3.095 1.410 ;
        RECT  2.705 1.150 2.935 1.310 ;
        RECT  2.545 0.425 2.705 1.310 ;
        RECT  1.645 0.425 2.545 0.585 ;
        RECT  1.385 0.385 1.645 0.635 ;
        RECT  0.720 0.475 1.385 0.635 ;
        RECT  0.560 0.475 0.720 1.580 ;
        RECT  0.430 1.205 0.560 1.580 ;
        END
        AntennaGateArea 0.2912 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 1.240 1.555 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.615 1.180 4.000 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.100 0.130 ;
        RECT  3.715 -0.130 3.975 0.980 ;
        RECT  0.835 -0.130 3.715 0.130 ;
        RECT  0.235 -0.130 0.835 0.285 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 1.870 3.975 3.000 ;
        RECT  1.290 2.740 3.715 3.000 ;
        RECT  0.690 2.165 1.290 3.000 ;
        RECT  0.000 2.740 0.690 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.275 0.370 3.435 2.360 ;
        RECT  2.885 0.370 3.275 0.970 ;
        RECT  3.175 1.760 3.275 2.360 ;
        RECT  2.025 1.930 2.365 2.190 ;
        RECT  1.635 2.400 2.155 2.560 ;
        RECT  1.865 0.815 2.025 2.190 ;
        RECT  1.235 0.815 1.865 0.975 ;
        RECT  1.475 1.760 1.635 2.560 ;
        RECT  0.250 1.760 1.475 1.920 ;
        RECT  0.250 0.765 0.335 1.025 ;
        RECT  0.090 0.765 0.250 1.920 ;
    END
END MXI2X2MTH

MACRO MXI2X3MTH
    CLASS CORE ;
    FOREIGN MXI2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.280 1.290 4.410 1.895 ;
        RECT  4.120 0.685 4.280 1.895 ;
        RECT  4.020 0.685 4.120 1.075 ;
        RECT  3.210 1.735 4.120 1.895 ;
        RECT  3.260 0.915 4.020 1.075 ;
        RECT  3.000 0.615 3.260 1.075 ;
        RECT  3.050 1.735 3.210 2.205 ;
        RECT  1.980 1.735 3.050 1.895 ;
        RECT  2.240 0.915 3.000 1.075 ;
        RECT  1.980 0.815 2.240 1.075 ;
        END
        AntennaDiffArea 1.34 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.200 1.390 1.580 ;
        END
        AntennaGateArea 0.4446 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 1.155 4.980 1.640 ;
        END
        AntennaGateArea 0.312 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.130 0.400 1.900 ;
        END
        AntennaGateArea 0.312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 0.255 ;
        RECT  1.670 -0.130 5.355 0.130 ;
        RECT  1.070 -0.130 1.670 0.265 ;
        RECT  0.000 -0.130 1.070 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.790 2.740 5.740 3.000 ;
        RECT  4.530 2.615 4.790 3.000 ;
        RECT  1.190 2.740 4.530 3.000 ;
        RECT  0.930 2.615 1.190 3.000 ;
        RECT  0.000 2.740 0.930 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.160 0.815 5.320 2.235 ;
        RECT  5.030 0.815 5.160 0.975 ;
        RECT  4.940 1.950 5.160 2.235 ;
        RECT  4.870 0.345 5.030 0.975 ;
        RECT  3.510 2.075 4.940 2.235 ;
        RECT  3.770 0.345 4.870 0.505 ;
        RECT  2.100 1.365 3.940 1.525 ;
        RECT  3.510 0.345 3.770 0.630 ;
        RECT  2.490 0.475 2.750 0.735 ;
        RECT  2.490 2.075 2.750 2.260 ;
        RECT  0.740 0.475 2.490 0.635 ;
        RECT  0.740 2.100 2.490 2.260 ;
        RECT  1.775 1.255 2.100 1.525 ;
        RECT  1.615 0.815 1.775 1.920 ;
        RECT  1.470 0.815 1.615 0.975 ;
        RECT  1.470 1.760 1.615 1.920 ;
        RECT  0.580 0.475 0.740 2.260 ;
    END
END MXI2X3MTH

MACRO MXI2X4MTH
    CLASS CORE ;
    FOREIGN MXI2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.795 0.775 4.975 1.990 ;
        RECT  3.455 0.775 4.795 0.955 ;
        RECT  4.265 1.700 4.795 1.990 ;
        RECT  3.565 1.700 4.265 1.880 ;
        RECT  3.305 1.700 3.565 2.365 ;
        RECT  3.195 0.355 3.455 0.955 ;
        RECT  2.540 1.700 3.305 1.880 ;
        RECT  2.520 0.775 3.195 0.955 ;
        RECT  2.280 1.700 2.540 1.975 ;
        RECT  2.360 0.685 2.520 0.955 ;
        RECT  2.175 0.685 2.360 0.845 ;
        END
        AntennaDiffArea 1.59 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.175 1.110 1.600 1.580 ;
        END
        AntennaGateArea 0.585 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.565 1.160 6.050 1.670 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.135 0.560 1.625 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 -0.130 6.150 0.130 ;
        RECT  5.765 -0.130 6.025 0.955 ;
        RECT  4.955 -0.130 5.765 0.130 ;
        RECT  4.695 -0.130 4.955 0.250 ;
        RECT  0.390 -0.130 4.695 0.130 ;
        RECT  0.130 -0.130 0.390 0.955 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 2.740 6.150 3.000 ;
        RECT  5.765 1.875 6.025 3.000 ;
        RECT  1.435 2.740 5.765 3.000 ;
        RECT  1.175 2.570 1.435 3.000 ;
        RECT  0.385 2.740 1.175 3.000 ;
        RECT  0.125 1.805 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.385 0.355 5.505 0.955 ;
        RECT  5.385 1.875 5.505 2.475 ;
        RECT  5.245 0.355 5.385 2.475 ;
        RECT  5.225 0.435 5.245 2.475 ;
        RECT  3.705 0.435 5.225 0.595 ;
        RECT  4.075 2.315 5.225 2.475 ;
        RECT  2.185 1.255 4.615 1.415 ;
        RECT  3.815 2.255 4.075 2.515 ;
        RECT  2.790 2.130 3.050 2.390 ;
        RECT  2.685 0.335 2.945 0.565 ;
        RECT  0.900 2.230 2.790 2.390 ;
        RECT  0.900 0.335 2.685 0.495 ;
        RECT  1.940 1.055 2.185 1.415 ;
        RECT  1.940 1.780 1.975 2.040 ;
        RECT  1.780 0.675 1.940 2.040 ;
        RECT  1.665 0.675 1.780 0.835 ;
        RECT  1.715 1.780 1.780 2.040 ;
        RECT  0.740 0.335 0.900 2.390 ;
        RECT  0.640 0.335 0.740 0.955 ;
        RECT  0.635 1.790 0.740 2.390 ;
    END
END MXI2X4MTH

MACRO MXI2X6MTH
    CLASS CORE ;
    FOREIGN MXI2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.720 0.800 6.990 1.990 ;
        RECT  4.870 0.800 6.720 1.070 ;
        RECT  6.660 1.635 6.720 1.990 ;
        RECT  4.995 1.720 6.660 1.990 ;
        RECT  4.735 1.720 4.995 2.420 ;
        RECT  4.610 0.425 4.870 1.070 ;
        RECT  3.710 1.720 4.735 1.990 ;
        RECT  3.850 0.800 4.610 1.070 ;
        RECT  3.590 0.765 3.850 1.070 ;
        END
        AntennaDiffArea 1.804 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.010 1.175 2.550 1.580 ;
        END
        AntennaGateArea 0.8801 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.525 1.210 8.145 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.250 1.065 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.965 -0.130 8.610 0.130 ;
        RECT  7.705 -0.130 7.965 0.615 ;
        RECT  0.900 -0.130 7.705 0.130 ;
        RECT  0.640 -0.130 0.900 0.615 ;
        RECT  0.000 -0.130 0.640 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.965 2.740 8.610 3.000 ;
        RECT  7.705 2.255 7.965 3.000 ;
        RECT  2.720 2.740 7.705 3.000 ;
        RECT  1.780 2.570 2.720 3.000 ;
        RECT  0.895 2.740 1.780 3.000 ;
        RECT  0.635 2.255 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.225 0.405 8.485 1.005 ;
        RECT  8.220 1.815 8.480 2.415 ;
        RECT  7.445 0.845 8.225 1.005 ;
        RECT  7.445 1.875 8.220 2.035 ;
        RECT  7.345 0.355 7.445 1.005 ;
        RECT  7.345 1.875 7.445 2.475 ;
        RECT  7.185 0.355 7.345 2.475 ;
        RECT  6.400 0.455 7.185 0.615 ;
        RECT  6.525 2.315 7.185 2.475 ;
        RECT  3.080 1.295 6.540 1.455 ;
        RECT  6.265 2.215 6.525 2.475 ;
        RECT  6.140 0.355 6.400 0.615 ;
        RECT  5.505 2.315 6.265 2.475 ;
        RECT  5.380 0.455 6.140 0.615 ;
        RECT  5.245 2.215 5.505 2.475 ;
        RECT  5.120 0.355 5.380 0.615 ;
        RECT  3.460 2.230 4.485 2.390 ;
        RECT  4.100 0.310 4.360 0.615 ;
        RECT  3.340 0.310 4.100 0.470 ;
        RECT  3.200 1.790 3.460 2.390 ;
        RECT  3.080 0.310 3.340 0.615 ;
        RECT  1.515 2.230 3.200 2.390 ;
        RECT  1.515 0.310 3.080 0.470 ;
        RECT  2.890 1.025 3.080 1.455 ;
        RECT  2.730 0.650 2.890 1.950 ;
        RECT  2.170 0.650 2.730 0.810 ;
        RECT  2.430 1.790 2.730 1.950 ;
        RECT  2.170 1.790 2.430 2.050 ;
        RECT  1.355 0.310 1.515 2.390 ;
        RECT  1.150 0.310 1.355 0.955 ;
        RECT  1.145 1.790 1.355 2.390 ;
        RECT  0.385 0.795 1.150 0.955 ;
        RECT  0.385 1.880 1.145 2.040 ;
        RECT  0.125 0.355 0.385 0.955 ;
        RECT  0.125 1.830 0.385 2.430 ;
    END
END MXI2X6MTH

MACRO MXI2X8MTH
    CLASS CORE ;
    FOREIGN MXI2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.380 0.785 8.680 2.025 ;
        RECT  6.020 0.785 8.380 1.095 ;
        RECT  6.110 1.695 8.380 2.025 ;
        RECT  5.850 1.695 6.110 2.400 ;
        RECT  5.760 0.395 6.020 1.095 ;
        RECT  3.805 1.695 5.850 2.025 ;
        RECT  3.960 0.785 5.760 1.095 ;
        RECT  3.750 0.710 3.960 1.095 ;
        END
        AntennaDiffArea 2.892 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.175 3.060 1.590 ;
        END
        AntennaGateArea 1.1739 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.345 1.225 10.305 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.230 1.580 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.595 -0.130 10.660 0.130 ;
        RECT  9.335 -0.130 9.595 0.620 ;
        RECT  1.405 -0.130 9.335 0.130 ;
        RECT  1.145 -0.130 1.405 0.615 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.960 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.595 2.740 10.660 3.000 ;
        RECT  9.335 2.255 9.595 3.000 ;
        RECT  3.555 2.740 9.335 3.000 ;
        RECT  3.295 2.550 3.555 3.000 ;
        RECT  2.455 2.740 3.295 3.000 ;
        RECT  2.195 2.550 2.455 3.000 ;
        RECT  1.405 2.740 2.195 3.000 ;
        RECT  1.145 2.255 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.905 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.855 0.380 10.115 0.980 ;
        RECT  9.855 1.855 10.115 2.455 ;
        RECT  9.075 0.820 9.855 0.980 ;
        RECT  9.075 1.855 9.855 2.015 ;
        RECT  8.915 0.365 9.075 2.515 ;
        RECT  8.865 0.365 8.915 0.980 ;
        RECT  8.815 2.255 8.915 2.515 ;
        RECT  6.270 0.405 8.865 0.565 ;
        RECT  7.645 2.355 8.815 2.515 ;
        RECT  3.540 1.315 8.200 1.475 ;
        RECT  7.385 2.255 7.645 2.515 ;
        RECT  6.620 2.355 7.385 2.515 ;
        RECT  6.360 2.255 6.620 2.515 ;
        RECT  5.340 2.255 5.600 2.515 ;
        RECT  5.230 0.310 5.490 0.565 ;
        RECT  4.575 2.255 5.340 2.415 ;
        RECT  4.470 0.310 5.230 0.470 ;
        RECT  4.315 2.255 4.575 2.515 ;
        RECT  4.210 0.310 4.470 0.565 ;
        RECT  3.895 2.255 4.315 2.415 ;
        RECT  1.920 0.310 4.210 0.470 ;
        RECT  3.735 2.210 3.895 2.415 ;
        RECT  1.920 2.210 3.735 2.370 ;
        RECT  3.380 0.650 3.540 1.475 ;
        RECT  2.260 0.650 3.380 0.810 ;
        RECT  2.755 1.770 3.015 2.030 ;
        RECT  2.260 1.770 2.755 1.930 ;
        RECT  2.100 0.650 2.260 1.930 ;
        RECT  1.760 0.310 1.920 2.370 ;
        RECT  1.655 0.310 1.760 0.970 ;
        RECT  1.655 1.770 1.760 2.370 ;
        RECT  0.895 0.810 1.655 0.970 ;
        RECT  0.895 1.770 1.655 1.930 ;
        RECT  0.635 0.370 0.895 0.970 ;
        RECT  0.635 1.770 0.895 2.425 ;
    END
END MXI2X8MTH

MACRO MXI2XLMTH
    CLASS CORE ;
    FOREIGN MXI2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.265 2.150 2.400 2.360 ;
        RECT  2.105 1.030 2.265 2.360 ;
        RECT  2.035 1.030 2.105 1.190 ;
        RECT  1.875 0.690 2.035 1.190 ;
        END
        AntennaDiffArea 0.352 ;
    END Y
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 0.310 1.735 0.470 ;
        RECT  1.475 0.310 1.635 0.635 ;
        RECT  0.720 0.475 1.475 0.635 ;
        RECT  0.560 0.475 0.720 1.610 ;
        RECT  0.430 1.245 0.560 1.610 ;
        END
        AntennaGateArea 0.1235 ;
    END S0
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.200 1.225 1.615 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.130 3.435 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.950 ;
        RECT  2.625 -0.130 3.305 0.390 ;
        RECT  1.295 -0.130 2.625 0.130 ;
        RECT  0.695 -0.130 1.295 0.285 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 2.740 3.690 3.000 ;
        RECT  3.305 1.800 3.565 3.000 ;
        RECT  2.965 2.490 3.305 3.000 ;
        RECT  0.905 2.740 2.965 3.000 ;
        RECT  0.745 2.135 0.905 3.000 ;
        RECT  0.000 2.740 0.745 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.775 0.740 2.995 0.900 ;
        RECT  2.775 1.770 2.835 2.030 ;
        RECT  2.615 0.740 2.775 2.030 ;
        RECT  2.395 0.740 2.615 0.900 ;
        RECT  1.765 1.370 1.925 2.345 ;
        RECT  1.245 2.185 1.765 2.345 ;
        RECT  1.425 0.815 1.585 2.005 ;
        RECT  1.255 0.815 1.425 0.975 ;
        RECT  1.085 1.795 1.245 2.345 ;
        RECT  0.250 1.795 1.085 1.955 ;
        RECT  0.250 0.765 0.335 1.025 ;
        RECT  0.090 0.765 0.250 1.955 ;
    END
END MXI2XLMTH

MACRO MXI3X1MTH
    CLASS CORE ;
    FOREIGN MXI3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.610 0.770 3.725 0.930 ;
        RECT  3.610 1.840 3.645 2.100 ;
        RECT  3.450 0.770 3.610 2.100 ;
        RECT  3.380 1.700 3.450 2.100 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 2.110 7.690 2.400 ;
        RECT  7.225 2.110 7.535 2.505 ;
        END
        AntennaGateArea 0.1612 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.095 0.515 2.400 ;
        END
        AntennaGateArea 0.1456 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.210 4.355 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.985 1.060 1.275 ;
        RECT  0.720 0.985 0.900 1.245 ;
        RECT  0.510 0.880 0.720 1.245 ;
        END
        AntennaGateArea 0.0884 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.880 3.180 1.520 ;
        RECT  2.675 1.205 2.970 1.520 ;
        END
        AntennaGateArea 0.0923 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.095 -0.130 7.790 0.130 ;
        RECT  6.835 -0.130 7.095 0.935 ;
        RECT  4.815 -0.130 6.835 0.130 ;
        RECT  4.215 -0.130 4.815 0.250 ;
        RECT  3.185 -0.130 4.215 0.130 ;
        RECT  2.585 -0.130 3.185 0.350 ;
        RECT  0.955 -0.130 2.585 0.130 ;
        RECT  0.695 -0.130 0.955 0.700 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 2.740 7.790 3.000 ;
        RECT  6.885 1.955 7.045 3.000 ;
        RECT  4.655 2.740 6.885 3.000 ;
        RECT  4.055 2.620 4.655 3.000 ;
        RECT  3.725 2.740 4.055 3.000 ;
        RECT  2.785 2.620 3.725 3.000 ;
        RECT  0.955 2.740 2.785 3.000 ;
        RECT  0.695 2.295 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.615 1.770 7.665 1.930 ;
        RECT  7.455 0.725 7.615 1.930 ;
        RECT  6.355 1.135 7.455 1.295 ;
        RECT  7.405 1.770 7.455 1.930 ;
        RECT  6.705 1.475 6.885 1.635 ;
        RECT  6.545 1.475 6.705 2.490 ;
        RECT  4.995 2.330 6.545 2.490 ;
        RECT  6.015 0.770 6.525 0.930 ;
        RECT  6.205 1.600 6.365 2.150 ;
        RECT  6.195 1.110 6.355 1.370 ;
        RECT  6.015 1.600 6.205 1.760 ;
        RECT  5.855 0.770 6.015 1.760 ;
        RECT  5.675 0.385 5.955 0.575 ;
        RECT  5.675 1.940 5.905 2.100 ;
        RECT  5.515 0.385 5.675 2.100 ;
        RECT  3.625 0.430 5.515 0.590 ;
        RECT  5.175 0.770 5.335 2.150 ;
        RECT  4.835 2.280 4.995 2.490 ;
        RECT  4.805 0.770 4.965 2.095 ;
        RECT  1.975 2.280 4.835 2.440 ;
        RECT  3.975 0.770 4.805 0.930 ;
        RECT  3.895 1.935 4.805 2.095 ;
        RECT  3.365 0.385 3.625 0.590 ;
        RECT  2.495 0.765 2.615 1.025 ;
        RECT  2.335 0.765 2.495 2.035 ;
        RECT  2.235 1.775 2.335 2.035 ;
        RECT  1.975 0.615 2.075 0.875 ;
        RECT  1.815 0.615 1.975 2.440 ;
        RECT  1.695 1.690 1.815 1.950 ;
        RECT  1.485 0.645 1.535 0.905 ;
        RECT  1.355 1.955 1.515 2.395 ;
        RECT  1.325 0.645 1.485 1.775 ;
        RECT  0.945 1.955 1.355 2.115 ;
        RECT  1.275 0.645 1.325 0.905 ;
        RECT  1.155 1.615 1.325 1.775 ;
        RECT  0.785 1.735 0.945 2.115 ;
        RECT  0.285 1.735 0.785 1.895 ;
        RECT  0.285 0.590 0.385 0.750 ;
        RECT  0.125 0.590 0.285 1.895 ;
    END
END MXI3X1MTH

MACRO MXI3X2MTH
    CLASS CORE ;
    FOREIGN MXI3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.300 0.360 8.510 2.310 ;
        RECT  8.225 0.360 8.300 0.960 ;
        RECT  8.225 1.710 8.300 2.310 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.495 1.110 6.870 1.580 ;
        END
        AntennaGateArea 0.2457 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.795 0.880 3.180 1.345 ;
        END
        AntennaGateArea 0.2054 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.700 1.185 4.000 1.665 ;
        END
        AntennaGateArea 0.0793 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.315 0.880 2.575 1.345 ;
        RECT  2.150 0.880 2.315 1.215 ;
        END
        AntennaGateArea 0.1261 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.965 0.355 1.845 ;
        END
        AntennaGateArea 0.1404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.600 -0.130 8.610 0.130 ;
        RECT  7.000 -0.130 7.600 0.250 ;
        RECT  4.410 -0.130 7.000 0.130 ;
        RECT  3.810 -0.130 4.410 0.250 ;
        RECT  2.505 -0.130 3.810 0.130 ;
        RECT  2.245 -0.130 2.505 0.700 ;
        RECT  0.385 -0.130 2.245 0.130 ;
        RECT  0.125 -0.130 0.385 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.975 2.740 8.610 3.000 ;
        RECT  7.815 1.685 7.975 3.000 ;
        RECT  7.715 1.685 7.815 1.945 ;
        RECT  7.260 2.620 7.815 3.000 ;
        RECT  4.275 2.740 7.260 3.000 ;
        RECT  3.675 2.620 4.275 3.000 ;
        RECT  2.475 2.740 3.675 3.000 ;
        RECT  2.315 2.205 2.475 3.000 ;
        RECT  0.725 2.740 2.315 3.000 ;
        RECT  0.125 2.615 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.045 1.165 8.095 1.425 ;
        RECT  7.885 0.430 8.045 1.425 ;
        RECT  5.410 0.430 7.885 0.590 ;
        RECT  7.055 2.250 7.625 2.410 ;
        RECT  7.210 0.770 7.480 0.930 ;
        RECT  7.210 1.810 7.365 2.070 ;
        RECT  7.050 0.770 7.210 2.070 ;
        RECT  6.895 2.250 7.055 2.560 ;
        RECT  6.715 1.910 7.050 2.070 ;
        RECT  4.615 2.400 6.895 2.560 ;
        RECT  6.555 1.910 6.715 2.220 ;
        RECT  5.785 2.060 6.555 2.220 ;
        RECT  6.310 0.770 6.480 0.930 ;
        RECT  6.310 1.720 6.375 1.880 ;
        RECT  6.150 0.770 6.310 1.880 ;
        RECT  6.115 1.180 6.150 1.880 ;
        RECT  5.930 1.180 6.115 1.440 ;
        RECT  5.750 0.770 5.970 0.930 ;
        RECT  5.750 1.960 5.785 2.220 ;
        RECT  5.590 0.770 5.750 2.220 ;
        RECT  5.325 0.430 5.410 1.560 ;
        RECT  5.250 0.430 5.325 2.110 ;
        RECT  5.165 1.400 5.250 2.110 ;
        RECT  5.065 1.850 5.165 2.110 ;
        RECT  4.765 0.525 4.950 0.785 ;
        RECT  4.765 1.900 4.815 2.060 ;
        RECT  4.605 0.525 4.765 2.060 ;
        RECT  4.455 2.280 4.615 2.560 ;
        RECT  4.555 1.900 4.605 2.060 ;
        RECT  2.815 2.280 4.455 2.440 ;
        RECT  4.340 1.370 4.410 1.630 ;
        RECT  4.180 0.790 4.340 2.075 ;
        RECT  3.860 0.790 4.180 0.950 ;
        RECT  3.455 1.915 4.180 2.075 ;
        RECT  3.700 0.690 3.860 0.950 ;
        RECT  3.360 0.540 3.520 1.685 ;
        RECT  2.995 0.540 3.360 0.700 ;
        RECT  3.155 1.525 3.360 1.685 ;
        RECT  2.995 1.525 3.155 2.075 ;
        RECT  2.135 1.525 2.995 1.685 ;
        RECT  2.655 1.865 2.815 2.440 ;
        RECT  2.135 1.865 2.655 2.025 ;
        RECT  1.975 1.395 2.135 1.685 ;
        RECT  1.975 1.865 2.135 2.335 ;
        RECT  1.765 1.395 1.975 1.555 ;
        RECT  1.305 2.175 1.975 2.335 ;
        RECT  1.695 0.715 1.955 1.115 ;
        RECT  1.635 1.735 1.795 1.995 ;
        RECT  1.605 1.295 1.765 1.555 ;
        RECT  1.425 0.955 1.695 1.115 ;
        RECT  1.425 1.735 1.635 1.895 ;
        RECT  1.265 0.955 1.425 1.895 ;
        RECT  1.085 0.605 1.415 0.765 ;
        RECT  1.085 2.075 1.305 2.335 ;
        RECT  0.925 0.605 1.085 2.335 ;
        RECT  0.585 0.640 0.745 2.095 ;
    END
END MXI3X2MTH

MACRO MXI3X4MTH
    CLASS CORE ;
    FOREIGN MXI3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.445 1.290 8.510 1.580 ;
        RECT  8.265 0.385 8.445 2.310 ;
        RECT  8.175 0.385 8.265 0.985 ;
        RECT  8.125 1.710 8.265 2.310 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.490 1.110 6.870 1.580 ;
        END
        AntennaGateArea 0.2574 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.815 0.880 3.180 1.335 ;
        END
        AntennaGateArea 0.2314 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 1.185 4.000 1.760 ;
        END
        AntennaGateArea 0.0871 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.315 0.880 2.575 1.335 ;
        RECT  2.150 0.880 2.315 1.170 ;
        END
        AntennaGateArea 0.1261 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.230 0.355 1.845 ;
        END
        AntennaGateArea 0.143 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 -0.130 9.020 0.130 ;
        RECT  8.635 -0.130 8.895 1.020 ;
        RECT  7.600 -0.130 8.635 0.130 ;
        RECT  7.000 -0.130 7.600 0.250 ;
        RECT  4.410 -0.130 7.000 0.130 ;
        RECT  3.810 -0.130 4.410 0.390 ;
        RECT  2.585 -0.130 3.810 0.130 ;
        RECT  2.325 -0.130 2.585 0.700 ;
        RECT  0.385 -0.130 2.325 0.130 ;
        RECT  0.125 -0.130 0.385 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 2.740 9.020 3.000 ;
        RECT  8.635 1.710 8.895 3.000 ;
        RECT  7.815 2.740 8.635 3.000 ;
        RECT  7.215 2.620 7.815 3.000 ;
        RECT  4.305 2.740 7.215 3.000 ;
        RECT  3.705 2.620 4.305 3.000 ;
        RECT  2.475 2.740 3.705 3.000 ;
        RECT  2.315 2.245 2.475 3.000 ;
        RECT  0.385 2.740 2.315 3.000 ;
        RECT  0.125 2.565 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.985 1.205 8.085 1.465 ;
        RECT  7.825 0.430 7.985 1.465 ;
        RECT  5.410 0.430 7.825 0.590 ;
        RECT  7.485 1.310 7.645 2.440 ;
        RECT  7.390 1.310 7.485 1.570 ;
        RECT  7.045 2.280 7.485 2.440 ;
        RECT  7.210 0.770 7.465 0.930 ;
        RECT  7.210 1.810 7.305 2.070 ;
        RECT  7.050 0.770 7.210 2.070 ;
        RECT  6.715 1.910 7.050 2.070 ;
        RECT  6.885 2.280 7.045 2.560 ;
        RECT  4.860 2.400 6.885 2.560 ;
        RECT  6.555 1.910 6.715 2.220 ;
        RECT  5.815 2.060 6.555 2.220 ;
        RECT  6.310 0.770 6.480 0.930 ;
        RECT  6.310 1.720 6.375 1.880 ;
        RECT  6.150 0.770 6.310 1.880 ;
        RECT  6.115 1.170 6.150 1.880 ;
        RECT  5.930 1.170 6.115 1.430 ;
        RECT  5.750 0.770 5.970 0.930 ;
        RECT  5.750 1.960 5.815 2.220 ;
        RECT  5.590 0.770 5.750 2.220 ;
        RECT  5.305 0.430 5.410 0.950 ;
        RECT  5.145 0.430 5.305 2.110 ;
        RECT  4.795 0.525 4.950 0.785 ;
        RECT  4.700 2.280 4.860 2.560 ;
        RECT  4.795 1.900 4.845 2.060 ;
        RECT  4.635 0.525 4.795 2.060 ;
        RECT  2.815 2.280 4.700 2.440 ;
        RECT  4.585 1.900 4.635 2.060 ;
        RECT  4.340 1.370 4.410 1.630 ;
        RECT  4.180 0.790 4.340 2.100 ;
        RECT  3.860 0.790 4.180 0.950 ;
        RECT  3.475 1.940 4.180 2.100 ;
        RECT  3.700 0.690 3.860 0.950 ;
        RECT  3.360 0.540 3.520 1.675 ;
        RECT  2.995 0.540 3.360 0.700 ;
        RECT  3.175 1.515 3.360 1.675 ;
        RECT  3.015 1.515 3.175 1.955 ;
        RECT  2.135 1.515 3.015 1.675 ;
        RECT  2.655 1.905 2.815 2.440 ;
        RECT  2.135 1.905 2.655 2.065 ;
        RECT  1.975 1.350 2.135 1.675 ;
        RECT  1.975 1.905 2.135 2.290 ;
        RECT  1.765 1.350 1.975 1.510 ;
        RECT  1.305 2.130 1.975 2.290 ;
        RECT  1.425 0.695 1.905 0.855 ;
        RECT  1.635 1.690 1.795 1.950 ;
        RECT  1.605 1.245 1.765 1.510 ;
        RECT  1.425 1.690 1.635 1.850 ;
        RECT  1.265 0.695 1.425 1.850 ;
        RECT  1.085 0.355 1.335 0.515 ;
        RECT  1.085 2.075 1.305 2.290 ;
        RECT  0.925 0.355 1.085 2.290 ;
        RECT  0.585 0.595 0.745 2.095 ;
    END
END MXI3X4MTH

MACRO MXI3X8MTH
    CLASS CORE ;
    FOREIGN MXI3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.310 0.420 9.660 2.385 ;
        RECT  9.120 0.745 9.310 2.125 ;
        RECT  8.615 0.745 9.120 1.095 ;
        RECT  8.640 1.775 9.120 2.125 ;
        RECT  8.290 1.775 8.640 2.385 ;
        RECT  8.385 0.420 8.615 1.095 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 0.880 6.870 1.495 ;
        RECT  6.495 1.235 6.660 1.495 ;
        END
        AntennaGateArea 0.2574 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.765 0.880 3.180 1.285 ;
        END
        AntennaGateArea 0.2314 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.725 1.185 4.105 1.670 ;
        END
        AntennaGateArea 0.0871 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.315 0.880 2.575 1.340 ;
        RECT  2.150 0.880 2.315 1.170 ;
        END
        AntennaGateArea 0.1261 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.230 0.405 1.845 ;
        END
        AntennaGateArea 0.143 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.085 -0.130 10.250 0.130 ;
        RECT  9.905 -0.130 10.085 1.020 ;
        RECT  9.105 -0.130 9.905 0.130 ;
        RECT  8.845 -0.130 9.105 0.565 ;
        RECT  8.055 -0.130 8.845 0.130 ;
        RECT  7.795 -0.130 8.055 0.250 ;
        RECT  7.055 -0.130 7.795 0.130 ;
        RECT  6.795 -0.130 7.055 0.250 ;
        RECT  4.390 -0.130 6.795 0.130 ;
        RECT  3.790 -0.130 4.390 0.385 ;
        RECT  2.585 -0.130 3.790 0.130 ;
        RECT  2.325 -0.130 2.585 0.700 ;
        RECT  0.385 -0.130 2.325 0.130 ;
        RECT  0.125 -0.130 0.385 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.085 2.740 10.250 3.000 ;
        RECT  9.905 1.710 10.085 3.000 ;
        RECT  9.105 2.740 9.905 3.000 ;
        RECT  8.845 2.305 9.105 3.000 ;
        RECT  8.025 2.740 8.845 3.000 ;
        RECT  7.425 2.620 8.025 3.000 ;
        RECT  4.390 2.740 7.425 3.000 ;
        RECT  3.790 2.620 4.390 3.000 ;
        RECT  2.475 2.740 3.790 3.000 ;
        RECT  2.315 2.245 2.475 3.000 ;
        RECT  0.385 2.740 2.315 3.000 ;
        RECT  0.125 2.620 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.195 1.315 8.765 1.475 ;
        RECT  8.035 0.430 8.195 1.475 ;
        RECT  5.410 0.430 8.035 0.590 ;
        RECT  7.695 1.410 7.855 2.440 ;
        RECT  7.550 1.410 7.695 1.570 ;
        RECT  7.255 2.280 7.695 2.440 ;
        RECT  7.210 0.770 7.605 0.930 ;
        RECT  7.390 1.310 7.550 1.570 ;
        RECT  7.210 1.810 7.515 2.070 ;
        RECT  7.095 2.280 7.255 2.560 ;
        RECT  7.050 0.770 7.210 2.070 ;
        RECT  4.795 2.400 7.095 2.560 ;
        RECT  6.925 1.910 7.050 2.070 ;
        RECT  6.765 1.910 6.925 2.220 ;
        RECT  5.950 2.060 6.765 2.220 ;
        RECT  6.310 1.720 6.585 1.880 ;
        RECT  6.310 0.795 6.480 0.955 ;
        RECT  6.150 0.795 6.310 1.880 ;
        RECT  5.930 1.180 6.150 1.440 ;
        RECT  5.750 0.770 5.970 0.930 ;
        RECT  5.750 1.960 5.950 2.220 ;
        RECT  5.590 0.770 5.750 2.220 ;
        RECT  5.230 0.430 5.410 2.110 ;
        RECT  4.795 0.525 4.955 2.060 ;
        RECT  4.690 0.525 4.795 0.785 ;
        RECT  4.670 1.900 4.795 2.060 ;
        RECT  4.635 2.280 4.795 2.560 ;
        RECT  2.815 2.280 4.635 2.440 ;
        RECT  4.450 1.360 4.540 1.620 ;
        RECT  4.290 0.690 4.450 2.015 ;
        RECT  3.700 0.690 4.290 0.950 ;
        RECT  3.475 1.855 4.290 2.015 ;
        RECT  3.360 0.540 3.520 1.625 ;
        RECT  2.995 0.540 3.360 0.700 ;
        RECT  3.175 1.465 3.360 1.625 ;
        RECT  3.015 1.465 3.175 1.945 ;
        RECT  2.135 1.520 3.015 1.680 ;
        RECT  2.655 1.905 2.815 2.440 ;
        RECT  2.135 1.905 2.655 2.065 ;
        RECT  1.975 1.350 2.135 1.680 ;
        RECT  1.975 1.905 2.135 2.290 ;
        RECT  1.765 1.350 1.975 1.510 ;
        RECT  1.305 2.130 1.975 2.290 ;
        RECT  1.645 0.470 1.905 0.970 ;
        RECT  1.635 1.690 1.795 1.950 ;
        RECT  1.605 1.250 1.765 1.510 ;
        RECT  1.425 0.810 1.645 0.970 ;
        RECT  1.425 1.690 1.635 1.850 ;
        RECT  1.265 0.810 1.425 1.850 ;
        RECT  1.085 0.470 1.335 0.630 ;
        RECT  1.085 2.075 1.305 2.290 ;
        RECT  0.925 0.470 1.085 2.290 ;
        RECT  0.585 0.640 0.745 2.095 ;
    END
END MXI3X8MTH

MACRO MXI3XLMTH
    CLASS CORE ;
    FOREIGN MXI3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.815 3.745 0.975 ;
        RECT  3.540 1.700 3.655 2.100 ;
        RECT  3.380 0.815 3.540 2.100 ;
        END
        AntennaDiffArea 0.226 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.245 2.110 7.690 2.505 ;
        END
        AntennaGateArea 0.1131 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.095 0.515 2.400 ;
        END
        AntennaGateArea 0.1066 ;
    END S0
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.025 1.260 4.420 1.725 ;
        END
        AntennaGateArea 0.0533 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.750 0.880 1.130 1.425 ;
        END
        AntennaGateArea 0.0533 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 1.145 3.180 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.095 -0.130 7.790 0.130 ;
        RECT  6.835 -0.130 7.095 1.015 ;
        RECT  4.785 -0.130 6.835 0.130 ;
        RECT  4.185 -0.130 4.785 0.250 ;
        RECT  3.165 -0.130 4.185 0.130 ;
        RECT  2.565 -0.130 3.165 0.350 ;
        RECT  0.955 -0.130 2.565 0.130 ;
        RECT  0.695 -0.130 0.955 0.700 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.045 2.740 7.790 3.000 ;
        RECT  6.885 1.875 7.045 3.000 ;
        RECT  4.705 2.740 6.885 3.000 ;
        RECT  4.105 2.620 4.705 3.000 ;
        RECT  3.595 2.740 4.105 3.000 ;
        RECT  2.995 2.620 3.595 3.000 ;
        RECT  0.955 2.740 2.995 3.000 ;
        RECT  0.695 2.295 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.405 0.765 7.665 1.930 ;
        RECT  6.345 1.195 7.405 1.355 ;
        RECT  6.705 1.535 6.885 1.695 ;
        RECT  6.545 1.535 6.705 2.520 ;
        RECT  5.130 2.360 6.545 2.520 ;
        RECT  6.005 0.815 6.515 0.975 ;
        RECT  6.205 1.600 6.365 2.115 ;
        RECT  6.185 1.160 6.345 1.420 ;
        RECT  6.005 1.600 6.205 1.760 ;
        RECT  5.845 0.815 6.005 1.760 ;
        RECT  5.665 0.430 5.945 0.635 ;
        RECT  5.665 1.940 5.845 2.100 ;
        RECT  5.505 0.430 5.665 2.100 ;
        RECT  3.355 0.430 5.505 0.590 ;
        RECT  5.165 0.770 5.325 2.100 ;
        RECT  5.015 1.940 5.165 2.100 ;
        RECT  4.970 2.280 5.130 2.520 ;
        RECT  4.835 1.485 4.985 1.745 ;
        RECT  2.055 2.280 4.970 2.440 ;
        RECT  4.675 0.820 4.835 2.065 ;
        RECT  3.995 0.820 4.675 0.980 ;
        RECT  3.955 1.905 4.675 2.065 ;
        RECT  2.565 0.635 2.675 0.895 ;
        RECT  2.565 1.785 2.675 2.045 ;
        RECT  2.405 0.635 2.565 2.045 ;
        RECT  1.895 0.635 2.055 2.440 ;
        RECT  1.525 1.955 1.685 2.355 ;
        RECT  1.375 0.635 1.535 1.775 ;
        RECT  0.945 1.955 1.525 2.115 ;
        RECT  1.325 0.635 1.375 0.895 ;
        RECT  1.275 1.615 1.375 1.775 ;
        RECT  0.785 1.735 0.945 2.115 ;
        RECT  0.385 1.735 0.785 1.895 ;
        RECT  0.125 0.635 0.385 1.895 ;
    END
END MXI3XLMTH

MACRO MXI4X1MTH
    CLASS CORE ;
    FOREIGN MXI4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.325 0.750 10.560 2.085 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 1.210 8.920 1.580 ;
        RECT  8.330 1.210 8.710 1.510 ;
        END
        AntennaGateArea 0.1612 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.480 0.880 3.590 1.270 ;
        RECT  3.380 0.880 3.480 1.430 ;
        RECT  3.290 1.080 3.380 1.430 ;
        END
        AntennaGateArea 0.2626 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 0.765 4.000 1.315 ;
        END
        AntennaGateArea 0.0923 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.780 0.880 6.050 1.460 ;
        RECT  5.630 1.200 5.780 1.460 ;
        END
        AntennaGateArea 0.0923 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 0.880 2.770 1.395 ;
        END
        AntennaGateArea 0.0923 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.120 0.395 1.580 ;
        END
        AntennaGateArea 0.0923 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.380 -0.130 10.660 0.130 ;
        RECT  9.780 -0.130 10.380 0.400 ;
        RECT  6.030 -0.130 9.780 0.130 ;
        RECT  5.770 -0.130 6.030 0.700 ;
        RECT  3.810 -0.130 5.770 0.130 ;
        RECT  3.550 -0.130 3.810 0.585 ;
        RECT  2.650 -0.130 3.550 0.130 ;
        RECT  2.390 -0.130 2.650 0.700 ;
        RECT  0.725 -0.130 2.390 0.130 ;
        RECT  0.125 -0.130 0.725 0.455 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 2.740 10.660 3.000 ;
        RECT  9.820 2.555 10.320 3.000 ;
        RECT  3.480 2.740 9.820 3.000 ;
        RECT  3.220 2.295 3.480 3.000 ;
        RECT  2.645 2.740 3.220 3.000 ;
        RECT  2.385 2.295 2.645 3.000 ;
        RECT  0.725 2.740 2.385 3.000 ;
        RECT  0.125 2.475 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.985 0.785 10.145 1.395 ;
        RECT  9.600 0.785 9.985 0.945 ;
        RECT  9.480 1.175 9.640 2.560 ;
        RECT  9.440 0.365 9.600 0.945 ;
        RECT  9.440 1.175 9.480 1.435 ;
        RECT  3.820 2.400 9.480 2.560 ;
        RECT  7.240 0.365 9.440 0.525 ;
        RECT  9.260 1.695 9.300 1.955 ;
        RECT  9.100 0.800 9.260 2.220 ;
        RECT  9.000 0.800 9.100 0.960 ;
        RECT  7.750 2.060 9.100 2.220 ;
        RECT  8.090 1.720 8.325 1.880 ;
        RECT  8.090 0.800 8.170 0.960 ;
        RECT  7.930 0.800 8.090 1.880 ;
        RECT  7.880 0.800 7.930 1.430 ;
        RECT  7.760 1.170 7.880 1.430 ;
        RECT  7.580 1.785 7.750 2.220 ;
        RECT  7.580 0.705 7.610 0.965 ;
        RECT  7.420 0.705 7.580 2.220 ;
        RECT  7.080 0.365 7.240 2.025 ;
        RECT  6.910 0.565 7.080 0.825 ;
        RECT  6.570 0.560 6.730 2.025 ;
        RECT  6.370 0.560 6.570 0.955 ;
        RECT  6.230 1.185 6.390 2.220 ;
        RECT  5.090 2.060 6.230 2.220 ;
        RECT  5.430 1.720 5.680 1.880 ;
        RECT  5.270 0.540 5.430 1.880 ;
        RECT  4.930 0.615 5.090 2.220 ;
        RECT  4.700 0.615 4.930 0.775 ;
        RECT  4.590 0.975 4.750 1.995 ;
        RECT  4.340 0.975 4.590 1.135 ;
        RECT  4.000 1.835 4.590 1.995 ;
        RECT  4.250 1.345 4.410 1.655 ;
        RECT  4.180 0.605 4.340 1.135 ;
        RECT  3.820 1.495 4.250 1.655 ;
        RECT  3.660 1.495 3.820 1.770 ;
        RECT  3.660 1.950 3.820 2.560 ;
        RECT  3.110 1.610 3.660 1.770 ;
        RECT  2.150 1.950 3.660 2.110 ;
        RECT  3.110 0.640 3.170 0.900 ;
        RECT  2.950 0.640 3.110 1.770 ;
        RECT  2.150 1.610 2.950 1.770 ;
        RECT  1.990 1.345 2.150 1.770 ;
        RECT  1.990 1.950 2.150 2.395 ;
        RECT  1.595 1.345 1.990 1.505 ;
        RECT  1.320 2.215 1.990 2.395 ;
        RECT  1.795 0.625 1.895 0.885 ;
        RECT  1.650 1.685 1.810 2.025 ;
        RECT  1.635 0.625 1.795 1.165 ;
        RECT  1.415 1.685 1.650 1.845 ;
        RECT  1.415 1.005 1.635 1.165 ;
        RECT  1.255 1.005 1.415 1.845 ;
        RECT  1.075 0.665 1.325 0.825 ;
        RECT  1.075 2.025 1.320 2.395 ;
        RECT  0.915 0.665 1.075 2.395 ;
        RECT  0.575 0.765 0.735 2.145 ;
    END
END MXI4X1MTH

MACRO MXI4X2MTH
    CLASS CORE ;
    FOREIGN MXI4X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.275 0.345 10.565 2.330 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.870 8.920 1.370 ;
        RECT  8.405 1.110 8.710 1.370 ;
        END
        AntennaGateArea 0.2327 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.880 3.590 1.400 ;
        RECT  2.985 1.240 3.380 1.400 ;
        END
        AntennaGateArea 0.4082 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 0.880 4.025 1.430 ;
        END
        AntennaGateArea 0.1261 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.815 0.880 6.155 1.540 ;
        END
        AntennaGateArea 0.1495 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.305 0.880 2.465 1.395 ;
        RECT  2.150 0.880 2.305 1.170 ;
        END
        AntennaGateArea 0.1248 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.875 0.395 1.750 ;
        END
        AntennaGateArea 0.1482 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.975 -0.130 10.660 0.130 ;
        RECT  9.815 -0.130 9.975 0.615 ;
        RECT  6.325 -0.130 9.815 0.130 ;
        RECT  6.065 -0.130 6.325 0.700 ;
        RECT  3.865 -0.130 6.065 0.130 ;
        RECT  3.605 -0.130 3.865 0.700 ;
        RECT  2.625 -0.130 3.605 0.130 ;
        RECT  2.365 -0.130 2.625 0.700 ;
        RECT  0.000 -0.130 2.365 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.025 2.740 10.660 3.000 ;
        RECT  9.765 1.855 10.025 3.000 ;
        RECT  3.715 2.740 9.765 3.000 ;
        RECT  3.455 2.295 3.715 3.000 ;
        RECT  2.625 2.740 3.455 3.000 ;
        RECT  2.365 2.295 2.625 3.000 ;
        RECT  0.725 2.740 2.365 3.000 ;
        RECT  0.125 2.565 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.935 0.795 10.095 1.395 ;
        RECT  9.635 0.795 9.935 0.955 ;
        RECT  9.475 0.365 9.635 0.955 ;
        RECT  9.295 1.750 9.485 2.220 ;
        RECT  7.375 0.365 9.475 0.525 ;
        RECT  9.135 0.750 9.295 2.220 ;
        RECT  4.055 2.400 9.225 2.560 ;
        RECT  7.885 2.060 9.135 2.220 ;
        RECT  8.225 1.720 8.445 1.880 ;
        RECT  8.225 0.710 8.405 0.870 ;
        RECT  8.065 0.710 8.225 1.880 ;
        RECT  7.895 1.170 8.065 1.430 ;
        RECT  7.715 1.865 7.885 2.220 ;
        RECT  7.715 0.705 7.845 0.965 ;
        RECT  7.555 0.705 7.715 2.220 ;
        RECT  7.145 0.365 7.375 2.025 ;
        RECT  6.705 0.565 6.865 2.025 ;
        RECT  6.585 0.565 6.705 0.825 ;
        RECT  6.365 1.335 6.525 2.220 ;
        RECT  5.295 2.060 6.365 2.220 ;
        RECT  5.635 1.720 5.885 1.880 ;
        RECT  5.635 0.540 5.805 0.700 ;
        RECT  5.475 0.540 5.635 1.880 ;
        RECT  5.035 0.485 5.295 2.220 ;
        RECT  4.685 0.725 4.845 2.165 ;
        RECT  4.205 0.725 4.685 0.985 ;
        RECT  4.235 2.005 4.685 2.165 ;
        RECT  4.345 1.255 4.505 1.775 ;
        RECT  2.805 1.615 4.345 1.775 ;
        RECT  3.895 1.955 4.055 2.560 ;
        RECT  2.125 1.955 3.895 2.115 ;
        RECT  2.955 0.500 3.115 1.040 ;
        RECT  2.805 0.880 2.955 1.040 ;
        RECT  2.645 0.880 2.805 1.775 ;
        RECT  2.125 1.615 2.645 1.775 ;
        RECT  1.965 1.350 2.125 1.775 ;
        RECT  1.965 1.955 2.125 2.310 ;
        RECT  1.595 1.350 1.965 1.510 ;
        RECT  1.295 2.130 1.965 2.310 ;
        RECT  1.755 0.535 1.915 1.170 ;
        RECT  1.625 1.690 1.785 1.950 ;
        RECT  1.415 1.010 1.755 1.170 ;
        RECT  1.415 1.690 1.625 1.850 ;
        RECT  1.075 0.570 1.455 0.830 ;
        RECT  1.255 1.010 1.415 1.850 ;
        RECT  1.075 2.055 1.295 2.310 ;
        RECT  0.915 0.570 1.075 2.310 ;
        RECT  0.575 0.730 0.735 2.050 ;
    END
END MXI4X2MTH

MACRO MXI4X4MTH
    CLASS CORE ;
    FOREIGN MXI4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 1.275 10.970 1.580 ;
        RECT  10.635 0.345 10.845 2.285 ;
        RECT  10.585 1.685 10.635 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 0.870 9.000 1.455 ;
        RECT  8.605 1.160 8.710 1.455 ;
        END
        AntennaGateArea 0.26 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.335 0.880 3.590 1.430 ;
        RECT  3.215 1.170 3.335 1.430 ;
        END
        AntennaGateArea 0.5005 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.880 4.175 1.395 ;
        END
        AntennaGateArea 0.1261 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.295 0.880 6.460 1.170 ;
        RECT  6.065 0.880 6.295 1.460 ;
        END
        AntennaGateArea 0.1755 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.305 0.880 2.550 1.395 ;
        RECT  2.150 0.880 2.305 1.170 ;
        END
        AntennaGateArea 0.1261 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.120 0.375 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 -0.130 11.480 0.130 ;
        RECT  11.095 -0.130 11.355 0.955 ;
        RECT  10.360 -0.130 11.095 0.130 ;
        RECT  10.125 -0.130 10.360 0.615 ;
        RECT  6.445 -0.130 10.125 0.130 ;
        RECT  6.185 -0.130 6.445 0.695 ;
        RECT  4.015 -0.130 6.185 0.130 ;
        RECT  3.755 -0.130 4.015 0.700 ;
        RECT  2.695 -0.130 3.755 0.130 ;
        RECT  2.435 -0.130 2.695 0.700 ;
        RECT  0.000 -0.130 2.435 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 2.740 11.480 3.000 ;
        RECT  11.095 1.865 11.355 3.000 ;
        RECT  10.335 2.740 11.095 3.000 ;
        RECT  10.075 1.890 10.335 3.000 ;
        RECT  3.865 2.740 10.075 3.000 ;
        RECT  3.605 2.295 3.865 3.000 ;
        RECT  2.695 2.740 3.605 3.000 ;
        RECT  2.435 2.295 2.695 3.000 ;
        RECT  0.000 2.740 2.435 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.290 0.795 10.450 1.465 ;
        RECT  9.945 0.795 10.290 0.955 ;
        RECT  9.785 0.340 9.945 0.955 ;
        RECT  9.605 1.825 9.825 2.220 ;
        RECT  7.435 0.340 9.785 0.500 ;
        RECT  9.445 0.705 9.605 2.220 ;
        RECT  4.205 2.400 9.565 2.560 ;
        RECT  9.345 0.705 9.445 0.865 ;
        RECT  7.915 2.060 9.445 2.220 ;
        RECT  8.395 1.720 8.645 1.880 ;
        RECT  8.395 0.720 8.520 0.980 ;
        RECT  8.235 0.720 8.395 1.880 ;
        RECT  8.095 1.195 8.235 1.455 ;
        RECT  7.915 0.705 8.010 0.965 ;
        RECT  7.755 0.705 7.915 2.220 ;
        RECT  7.435 1.765 7.575 2.025 ;
        RECT  7.275 0.340 7.435 2.025 ;
        RECT  6.935 0.660 7.095 2.025 ;
        RECT  6.705 0.660 6.935 0.920 ;
        RECT  6.905 1.765 6.935 2.025 ;
        RECT  6.655 1.365 6.755 1.525 ;
        RECT  6.495 1.365 6.655 2.220 ;
        RECT  5.445 2.060 6.495 2.220 ;
        RECT  5.785 1.720 6.065 1.880 ;
        RECT  5.785 0.540 5.925 0.700 ;
        RECT  5.625 0.540 5.785 1.880 ;
        RECT  5.365 1.805 5.445 2.220 ;
        RECT  5.205 0.485 5.365 2.220 ;
        RECT  4.835 0.685 4.995 2.165 ;
        RECT  4.355 0.685 4.835 0.945 ;
        RECT  4.385 2.005 4.835 2.165 ;
        RECT  4.495 1.315 4.655 1.770 ;
        RECT  3.035 1.610 4.495 1.770 ;
        RECT  4.045 1.955 4.205 2.560 ;
        RECT  2.125 1.955 4.045 2.115 ;
        RECT  3.035 0.600 3.155 0.860 ;
        RECT  2.875 0.600 3.035 1.770 ;
        RECT  2.125 1.610 2.875 1.770 ;
        RECT  1.965 1.350 2.125 1.770 ;
        RECT  1.965 1.955 2.125 2.310 ;
        RECT  1.745 1.350 1.965 1.510 ;
        RECT  1.295 2.130 1.965 2.310 ;
        RECT  1.705 0.535 1.865 1.170 ;
        RECT  1.625 1.690 1.785 1.950 ;
        RECT  1.415 1.010 1.705 1.170 ;
        RECT  1.415 1.690 1.625 1.850 ;
        RECT  1.255 1.010 1.415 1.850 ;
        RECT  1.075 0.570 1.325 0.830 ;
        RECT  1.075 2.055 1.295 2.310 ;
        RECT  0.915 0.570 1.075 2.310 ;
        RECT  0.575 0.765 0.735 1.965 ;
    END
END MXI4X4MTH

MACRO MXI4X8MTH
    CLASS CORE ;
    FOREIGN MXI4X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.360 0.380 11.710 2.360 ;
        RECT  10.765 1.205 11.360 1.555 ;
        RECT  10.465 0.380 10.765 2.350 ;
        RECT  10.385 0.380 10.465 0.980 ;
        RECT  10.385 1.750 10.465 2.350 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.635 0.880 8.920 1.470 ;
        RECT  8.565 1.190 8.635 1.470 ;
        END
        AntennaGateArea 0.26 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.880 3.590 1.420 ;
        RECT  3.215 1.160 3.380 1.420 ;
        END
        AntennaGateArea 0.5005 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.880 4.175 1.430 ;
        END
        AntennaGateArea 0.1261 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.260 0.880 6.460 1.170 ;
        RECT  6.055 0.880 6.260 1.460 ;
        END
        AntennaGateArea 0.1755 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.305 0.880 2.510 1.395 ;
        RECT  2.150 0.880 2.305 1.175 ;
        END
        AntennaGateArea 0.1261 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.120 0.375 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 -0.130 12.300 0.130 ;
        RECT  11.915 -0.130 12.175 0.980 ;
        RECT  11.105 -0.130 11.915 0.130 ;
        RECT  10.945 -0.130 11.105 0.980 ;
        RECT  10.055 -0.130 10.945 0.130 ;
        RECT  9.795 -0.130 10.055 0.250 ;
        RECT  6.445 -0.130 9.795 0.130 ;
        RECT  6.185 -0.130 6.445 0.695 ;
        RECT  3.995 -0.130 6.185 0.130 ;
        RECT  3.735 -0.130 3.995 0.585 ;
        RECT  2.695 -0.130 3.735 0.130 ;
        RECT  2.435 -0.130 2.695 0.700 ;
        RECT  0.000 -0.130 2.435 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.175 2.740 12.300 3.000 ;
        RECT  11.915 1.860 12.175 3.000 ;
        RECT  11.105 2.740 11.915 3.000 ;
        RECT  10.945 1.865 11.105 3.000 ;
        RECT  3.865 2.740 10.945 3.000 ;
        RECT  3.605 2.295 3.865 3.000 ;
        RECT  2.695 2.740 3.605 3.000 ;
        RECT  2.435 2.295 2.695 3.000 ;
        RECT  0.000 2.740 2.435 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.205 1.205 10.285 1.465 ;
        RECT  10.045 0.430 10.205 1.465 ;
        RECT  9.040 0.430 10.045 0.590 ;
        RECT  9.400 1.695 9.685 1.955 ;
        RECT  9.400 0.795 9.500 0.955 ;
        RECT  4.205 2.400 9.425 2.560 ;
        RECT  9.240 0.795 9.400 2.220 ;
        RECT  7.925 2.060 9.240 2.220 ;
        RECT  8.765 0.340 9.040 0.590 ;
        RECT  7.435 0.340 8.765 0.500 ;
        RECT  8.340 1.720 8.655 1.880 ;
        RECT  8.340 0.750 8.455 1.010 ;
        RECT  8.180 0.750 8.340 1.880 ;
        RECT  8.105 1.195 8.180 1.455 ;
        RECT  7.925 0.705 7.995 0.965 ;
        RECT  7.765 0.705 7.925 2.220 ;
        RECT  7.435 1.765 7.585 2.025 ;
        RECT  7.275 0.340 7.435 2.025 ;
        RECT  6.935 0.685 7.095 2.025 ;
        RECT  6.705 0.685 6.935 0.845 ;
        RECT  6.885 1.765 6.935 2.025 ;
        RECT  6.655 1.365 6.755 1.525 ;
        RECT  6.495 1.365 6.655 2.220 ;
        RECT  5.475 2.060 6.495 2.220 ;
        RECT  5.825 1.720 6.065 1.880 ;
        RECT  5.825 0.540 5.925 0.700 ;
        RECT  5.665 0.540 5.825 1.880 ;
        RECT  5.365 1.960 5.475 2.220 ;
        RECT  5.205 0.485 5.365 2.220 ;
        RECT  4.835 0.665 4.995 2.215 ;
        RECT  4.355 0.665 4.835 0.925 ;
        RECT  4.385 1.955 4.835 2.215 ;
        RECT  4.495 1.315 4.655 1.770 ;
        RECT  3.035 1.610 4.495 1.770 ;
        RECT  4.045 1.955 4.205 2.560 ;
        RECT  2.125 1.955 4.045 2.115 ;
        RECT  3.035 0.600 3.155 0.860 ;
        RECT  2.875 0.600 3.035 1.770 ;
        RECT  2.125 1.610 2.875 1.770 ;
        RECT  1.965 1.360 2.125 1.770 ;
        RECT  1.965 1.955 2.125 2.320 ;
        RECT  1.745 1.360 1.965 1.520 ;
        RECT  1.295 2.140 1.965 2.320 ;
        RECT  1.705 0.535 1.865 1.175 ;
        RECT  1.625 1.700 1.785 1.960 ;
        RECT  1.565 1.015 1.705 1.175 ;
        RECT  1.565 1.700 1.625 1.860 ;
        RECT  1.405 1.015 1.565 1.860 ;
        RECT  1.075 0.560 1.325 0.830 ;
        RECT  1.075 2.055 1.295 2.320 ;
        RECT  0.915 0.560 1.075 2.320 ;
        RECT  0.575 0.765 0.735 1.965 ;
    END
END MXI4X8MTH

MACRO MXI4XLMTH
    CLASS CORE ;
    FOREIGN MXI4XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.325 0.750 10.560 1.990 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN S1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 1.210 8.920 1.580 ;
        RECT  8.330 1.210 8.710 1.510 ;
        END
        AntennaGateArea 0.1131 ;
    END S1
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 0.880 3.590 1.270 ;
        RECT  3.380 0.880 3.450 1.430 ;
        RECT  3.290 1.080 3.380 1.430 ;
        END
        AntennaGateArea 0.1599 ;
    END S0
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 0.765 4.000 1.300 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.930 0.880 6.090 1.130 ;
        RECT  5.680 0.880 5.930 1.460 ;
        END
        AntennaGateArea 0.0624 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 0.880 2.770 1.395 ;
        END
        AntennaGateArea 0.0533 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.120 0.395 1.580 ;
        END
        AntennaGateArea 0.078 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.380 -0.130 10.660 0.130 ;
        RECT  9.780 -0.130 10.380 0.400 ;
        RECT  9.480 -0.130 9.780 0.130 ;
        RECT  8.540 -0.130 9.480 0.250 ;
        RECT  6.395 -0.130 8.540 0.130 ;
        RECT  5.455 -0.130 6.395 0.315 ;
        RECT  3.810 -0.130 5.455 0.130 ;
        RECT  3.550 -0.130 3.810 0.585 ;
        RECT  2.650 -0.130 3.550 0.130 ;
        RECT  2.390 -0.130 2.650 0.700 ;
        RECT  0.725 -0.130 2.390 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.320 2.740 10.660 3.000 ;
        RECT  9.820 2.375 10.320 3.000 ;
        RECT  3.450 2.740 9.820 3.000 ;
        RECT  3.190 2.295 3.450 3.000 ;
        RECT  2.590 2.740 3.190 3.000 ;
        RECT  2.330 2.295 2.590 3.000 ;
        RECT  0.725 2.740 2.330 3.000 ;
        RECT  0.125 2.245 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.955 0.785 10.115 1.445 ;
        RECT  9.600 0.785 9.955 0.945 ;
        RECT  9.480 1.205 9.640 2.560 ;
        RECT  9.440 0.460 9.600 0.945 ;
        RECT  9.440 1.205 9.480 1.465 ;
        RECT  3.790 2.400 9.480 2.560 ;
        RECT  8.320 0.460 9.440 0.620 ;
        RECT  9.260 1.695 9.300 2.220 ;
        RECT  9.100 0.800 9.260 2.220 ;
        RECT  9.000 0.800 9.100 0.960 ;
        RECT  7.750 2.060 9.100 2.220 ;
        RECT  8.090 1.720 8.325 1.880 ;
        RECT  8.065 0.365 8.320 0.620 ;
        RECT  8.090 0.800 8.230 0.960 ;
        RECT  7.930 0.800 8.090 1.880 ;
        RECT  7.180 0.365 8.065 0.525 ;
        RECT  7.760 1.170 7.930 1.430 ;
        RECT  7.580 1.715 7.750 2.220 ;
        RECT  7.580 0.705 7.670 0.965 ;
        RECT  7.420 0.705 7.580 2.220 ;
        RECT  7.020 0.365 7.180 1.975 ;
        RECT  6.940 0.365 7.020 0.825 ;
        RECT  6.620 0.970 6.780 1.930 ;
        RECT  6.530 0.970 6.620 1.130 ;
        RECT  6.450 1.670 6.620 1.930 ;
        RECT  6.370 0.565 6.530 1.130 ;
        RECT  6.270 1.310 6.440 1.470 ;
        RECT  6.110 1.310 6.270 2.220 ;
        RECT  5.090 2.060 6.110 2.220 ;
        RECT  5.430 1.720 5.710 1.880 ;
        RECT  5.430 0.565 5.490 0.825 ;
        RECT  5.270 0.565 5.430 1.880 ;
        RECT  4.930 0.615 5.090 2.220 ;
        RECT  4.700 0.615 4.930 0.775 ;
        RECT  4.590 0.975 4.750 1.980 ;
        RECT  4.340 0.975 4.590 1.135 ;
        RECT  3.970 1.820 4.590 1.980 ;
        RECT  4.250 1.315 4.410 1.640 ;
        RECT  4.180 0.605 4.340 1.135 ;
        RECT  3.790 1.480 4.250 1.640 ;
        RECT  3.630 1.480 3.790 1.770 ;
        RECT  3.630 1.950 3.790 2.560 ;
        RECT  3.110 1.610 3.630 1.770 ;
        RECT  2.150 1.950 3.630 2.110 ;
        RECT  3.110 0.625 3.170 0.885 ;
        RECT  2.950 0.625 3.110 1.770 ;
        RECT  2.150 1.610 2.950 1.770 ;
        RECT  1.990 1.355 2.150 1.770 ;
        RECT  1.990 1.950 2.150 2.315 ;
        RECT  1.595 1.355 1.990 1.515 ;
        RECT  1.355 2.135 1.990 2.315 ;
        RECT  1.635 0.625 1.895 1.175 ;
        RECT  1.415 1.695 1.810 1.955 ;
        RECT  1.415 1.015 1.635 1.175 ;
        RECT  1.255 1.015 1.415 1.955 ;
        RECT  1.075 2.135 1.355 2.425 ;
        RECT  1.075 0.670 1.325 0.830 ;
        RECT  0.915 0.670 1.075 2.425 ;
        RECT  0.575 0.765 0.735 1.945 ;
    END
END MXI4XLMTH

MACRO NAND2BX12MTH
    CLASS CORE ;
    FOREIGN NAND2BX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.740 0.435 8.070 2.310 ;
        RECT  2.850 0.435 7.740 0.805 ;
        RECT  7.555 1.535 7.740 2.310 ;
        RECT  7.160 1.535 7.555 2.500 ;
        RECT  2.250 1.960 7.160 2.500 ;
        END
        AntennaDiffArea 2.82 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.295 1.025 7.555 1.345 ;
        RECT  5.895 1.025 7.295 1.185 ;
        RECT  5.635 1.025 5.895 1.400 ;
        RECT  4.190 1.025 5.635 1.185 ;
        RECT  3.590 1.025 4.190 1.400 ;
        RECT  2.480 1.025 3.590 1.185 ;
        RECT  2.110 0.920 2.480 1.400 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.770 1.210 1.475 1.470 ;
        RECT  0.445 1.210 0.770 1.540 ;
        END
        AntennaGateArea 0.5304 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.810 -0.130 8.200 0.130 ;
        RECT  7.210 -0.130 7.810 0.255 ;
        RECT  5.750 -0.130 7.210 0.130 ;
        RECT  5.490 -0.130 5.750 0.255 ;
        RECT  4.020 -0.130 5.490 0.130 ;
        RECT  3.760 -0.130 4.020 0.255 ;
        RECT  2.255 -0.130 3.760 0.130 ;
        RECT  1.995 -0.130 2.255 0.735 ;
        RECT  1.140 -0.130 1.995 0.130 ;
        RECT  0.880 -0.130 1.140 0.640 ;
        RECT  0.000 -0.130 0.880 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.055 2.740 8.200 3.000 ;
        RECT  7.795 2.490 8.055 3.000 ;
        RECT  2.005 2.740 7.795 3.000 ;
        RECT  1.745 2.135 2.005 3.000 ;
        RECT  0.925 2.740 1.745 3.000 ;
        RECT  0.665 2.100 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.370 1.365 6.630 1.740 ;
        RECT  5.060 1.580 6.370 1.740 ;
        RECT  4.460 1.365 5.060 1.740 ;
        RECT  3.320 1.580 4.460 1.740 ;
        RECT  2.720 1.365 3.320 1.740 ;
        RECT  1.815 1.580 2.720 1.740 ;
        RECT  1.655 0.615 1.815 1.880 ;
        RECT  1.420 0.615 1.655 0.980 ;
        RECT  1.465 1.720 1.655 1.880 ;
        RECT  1.205 1.720 1.465 2.360 ;
        RECT  0.600 0.820 1.420 0.980 ;
        RECT  0.385 1.720 1.205 1.880 ;
        RECT  0.340 0.615 0.600 0.980 ;
        RECT  0.125 1.720 0.385 2.360 ;
    END
END NAND2BX12MTH

MACRO NAND2BX1MTH
    CLASS CORE ;
    FOREIGN NAND2BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 0.470 1.960 1.930 ;
        RECT  1.555 0.470 1.800 0.840 ;
        RECT  1.325 1.770 1.800 1.930 ;
        RECT  1.165 1.770 1.325 2.085 ;
        END
        AntennaDiffArea 0.36 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.820 1.225 1.250 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 0.880 0.720 1.240 ;
        RECT  0.460 0.880 0.645 1.550 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.955 -0.130 2.050 0.130 ;
        RECT  0.695 -0.130 0.955 0.640 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 2.740 2.050 3.000 ;
        RECT  1.655 2.110 1.915 3.000 ;
        RECT  1.375 2.740 1.655 3.000 ;
        RECT  1.115 2.570 1.375 3.000 ;
        RECT  0.825 2.740 1.115 3.000 ;
        RECT  0.225 2.195 0.825 3.000 ;
        RECT  0.000 2.740 0.225 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.405 1.095 1.620 1.590 ;
        RECT  0.985 1.430 1.405 1.590 ;
        RECT  0.825 1.430 0.985 1.895 ;
        RECT  0.250 1.735 0.825 1.895 ;
        RECT  0.250 0.490 0.335 0.750 ;
        RECT  0.090 0.490 0.250 1.895 ;
    END
END NAND2BX1MTH

MACRO NAND2BX2MTH
    CLASS CORE ;
    FOREIGN NAND2BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 0.470 1.950 2.260 ;
        RECT  1.535 0.470 1.790 0.760 ;
        RECT  1.385 2.100 1.790 2.260 ;
        RECT  1.125 2.100 1.385 2.360 ;
        END
        AntennaDiffArea 0.575 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 1.280 1.185 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.280 0.555 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.925 -0.130 2.050 0.130 ;
        RECT  0.665 -0.130 0.925 0.760 ;
        RECT  0.315 -0.130 0.665 0.360 ;
        RECT  0.000 -0.130 0.315 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 2.740 2.050 3.000 ;
        RECT  1.665 2.440 1.925 3.000 ;
        RECT  0.835 2.740 1.665 3.000 ;
        RECT  0.235 2.335 0.835 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.415 0.940 1.575 1.920 ;
        RECT  0.385 0.940 1.415 1.100 ;
        RECT  0.125 1.760 1.415 1.920 ;
        RECT  0.125 0.765 0.385 1.100 ;
    END
END NAND2BX2MTH

MACRO NAND2BX4MTH
    CLASS CORE ;
    FOREIGN NAND2BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 1.765 2.605 2.400 ;
        RECT  2.325 0.815 2.505 2.400 ;
        RECT  1.785 0.815 2.325 0.995 ;
        RECT  2.150 2.100 2.325 2.400 ;
        RECT  1.480 2.100 2.150 2.280 ;
        RECT  1.220 2.100 1.480 2.360 ;
        END
        AntennaDiffArea 0.938 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 1.135 2.945 1.395 ;
        RECT  2.685 0.475 2.845 1.395 ;
        RECT  1.240 0.475 2.685 0.635 ;
        RECT  1.080 0.475 1.240 1.480 ;
        RECT  0.920 0.880 1.080 1.480 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.090 0.400 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 -0.130 3.280 0.130 ;
        RECT  2.650 -0.130 2.910 0.250 ;
        RECT  1.130 -0.130 2.650 0.130 ;
        RECT  0.870 -0.130 1.130 0.295 ;
        RECT  0.000 -0.130 0.870 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.895 1.765 3.155 3.000 ;
        RECT  1.970 2.740 2.895 3.000 ;
        RECT  1.770 2.460 1.970 3.000 ;
        RECT  0.930 2.740 1.770 3.000 ;
        RECT  0.670 2.100 0.930 3.000 ;
        RECT  0.000 2.740 0.670 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.660 1.225 2.145 1.485 ;
        RECT  1.500 1.225 1.660 1.920 ;
        RECT  0.740 1.760 1.500 1.920 ;
        RECT  0.580 0.610 0.740 1.920 ;
        RECT  0.330 0.610 0.580 0.870 ;
        RECT  0.385 1.760 0.580 1.920 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END NAND2BX4MTH

MACRO NAND2BX8MTH
    CLASS CORE ;
    FOREIGN NAND2BX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.350 0.475 5.640 1.925 ;
        RECT  2.320 0.475 5.350 0.805 ;
        RECT  5.110 1.575 5.350 1.925 ;
        RECT  4.760 1.575 5.110 2.310 ;
        RECT  4.045 1.960 4.760 2.310 ;
        RECT  3.665 1.960 4.045 2.460 ;
        RECT  3.080 1.960 3.665 2.310 ;
        RECT  2.670 1.960 3.080 2.460 ;
        RECT  1.715 2.110 2.670 2.460 ;
        END
        AntennaDiffArea 1.882 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.940 1.025 5.170 1.395 ;
        RECT  3.655 1.025 4.940 1.185 ;
        RECT  3.055 1.025 3.655 1.400 ;
        RECT  1.990 1.025 3.055 1.185 ;
        RECT  1.440 1.025 1.990 1.540 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.195 0.805 1.540 ;
        END
        AntennaGateArea 0.3536 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.555 -0.130 5.740 0.130 ;
        RECT  4.955 -0.130 5.555 0.255 ;
        RECT  3.485 -0.130 4.955 0.130 ;
        RECT  3.225 -0.130 3.485 0.255 ;
        RECT  1.720 -0.130 3.225 0.130 ;
        RECT  1.460 -0.130 1.720 0.845 ;
        RECT  0.605 -0.130 1.460 0.130 ;
        RECT  0.345 -0.130 0.605 1.015 ;
        RECT  0.000 -0.130 0.345 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 2.105 5.615 3.000 ;
        RECT  4.525 2.740 5.355 3.000 ;
        RECT  4.265 2.490 4.525 3.000 ;
        RECT  1.470 2.740 4.265 3.000 ;
        RECT  1.210 2.135 1.470 3.000 ;
        RECT  0.390 2.740 1.210 3.000 ;
        RECT  0.130 1.790 0.390 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.925 1.365 4.525 1.740 ;
        RECT  2.785 1.580 3.925 1.740 ;
        RECT  2.345 1.365 2.785 1.740 ;
        RECT  2.185 1.365 2.345 1.880 ;
        RECT  1.145 1.720 2.185 1.880 ;
        RECT  0.985 0.615 1.145 1.880 ;
        RECT  0.885 0.615 0.985 0.875 ;
        RECT  0.930 1.720 0.985 1.880 ;
        RECT  0.670 1.720 0.930 2.360 ;
    END
END NAND2BX8MTH

MACRO NAND2BXLMTH
    CLASS CORE ;
    FOREIGN NAND2BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 0.470 1.960 1.925 ;
        RECT  1.585 0.470 1.800 0.805 ;
        RECT  1.440 1.765 1.800 1.925 ;
        RECT  1.180 1.765 1.440 2.025 ;
        END
        AntennaDiffArea 0.241 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.820 1.225 1.245 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 0.880 0.720 1.240 ;
        RECT  0.445 0.880 0.645 1.465 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 -0.130 2.050 0.130 ;
        RECT  0.955 -0.130 1.310 0.300 ;
        RECT  0.695 -0.130 0.955 0.640 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 2.740 2.050 3.000 ;
        RECT  1.325 2.480 1.925 3.000 ;
        RECT  1.145 2.740 1.325 3.000 ;
        RECT  0.205 2.480 1.145 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.405 1.095 1.620 1.585 ;
        RECT  0.985 1.425 1.405 1.585 ;
        RECT  0.825 1.425 0.985 1.915 ;
        RECT  0.250 1.755 0.825 1.915 ;
        RECT  0.250 0.475 0.335 0.735 ;
        RECT  0.090 0.475 0.250 1.915 ;
    END
END NAND2BXLMTH

MACRO NAND2X12MTH
    CLASS CORE ;
    FOREIGN NAND2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.130 0.430 6.430 2.440 ;
        RECT  1.205 0.430 6.130 0.790 ;
        RECT  5.615 1.495 6.130 2.440 ;
        RECT  4.655 1.865 5.615 2.440 ;
        RECT  3.865 1.865 4.655 2.125 ;
        RECT  3.605 1.865 3.865 2.475 ;
        RECT  2.905 1.865 3.605 2.125 ;
        RECT  2.645 1.865 2.905 2.465 ;
        RECT  1.925 1.865 2.645 2.125 ;
        RECT  1.665 1.865 1.925 2.465 ;
        RECT  0.905 1.865 1.665 2.125 ;
        RECT  0.645 1.865 0.905 2.465 ;
        END
        AntennaDiffArea 2.816 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.785 1.010 5.945 1.270 ;
        RECT  4.205 1.010 5.785 1.170 ;
        RECT  3.945 1.010 4.205 1.345 ;
        RECT  2.535 1.010 3.945 1.170 ;
        RECT  2.190 1.010 2.535 1.345 ;
        RECT  1.935 0.980 2.190 1.345 ;
        RECT  1.110 0.980 1.935 1.140 ;
        RECT  0.785 0.980 1.110 1.580 ;
        RECT  0.305 1.160 0.785 1.580 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.785 1.350 5.045 1.685 ;
        RECT  3.285 1.525 4.785 1.685 ;
        RECT  3.025 1.350 3.285 1.685 ;
        RECT  1.595 1.525 3.025 1.685 ;
        RECT  1.290 1.330 1.595 1.685 ;
        END
        AntennaGateArea 1.2324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.105 -0.130 6.560 0.130 ;
        RECT  5.505 -0.130 6.105 0.250 ;
        RECT  4.045 -0.130 5.505 0.130 ;
        RECT  3.785 -0.130 4.045 0.250 ;
        RECT  2.325 -0.130 3.785 0.130 ;
        RECT  2.065 -0.130 2.325 0.250 ;
        RECT  0.605 -0.130 2.065 0.130 ;
        RECT  0.345 -0.130 0.605 0.980 ;
        RECT  0.000 -0.130 0.345 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.425 2.740 6.560 3.000 ;
        RECT  6.165 2.620 6.425 3.000 ;
        RECT  4.385 2.740 6.165 3.000 ;
        RECT  4.125 2.305 4.385 3.000 ;
        RECT  1.415 2.740 4.125 3.000 ;
        RECT  1.155 2.305 1.415 3.000 ;
        RECT  0.385 2.740 1.155 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND2X12MTH

MACRO NAND2X1MTH
    CLASS CORE ;
    FOREIGN NAND2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.045 0.735 1.365 0.995 ;
        RECT  1.045 1.700 1.130 1.990 ;
        RECT  0.885 0.735 1.045 1.990 ;
        RECT  0.675 1.710 0.885 1.990 ;
        END
        AntennaDiffArea 0.36 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 0.705 1.465 ;
        RECT  0.100 1.205 0.310 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.250 1.540 1.990 ;
        RECT  1.225 1.250 1.330 1.510 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.165 -0.130 1.640 0.130 ;
        RECT  0.485 -0.130 1.165 0.300 ;
        RECT  0.225 -0.130 0.485 1.025 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 2.740 1.640 3.000 ;
        RECT  1.245 2.170 1.505 3.000 ;
        RECT  0.935 2.740 1.245 3.000 ;
        RECT  0.675 2.570 0.935 3.000 ;
        RECT  0.385 2.740 0.675 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND2X1MTH

MACRO NAND2X2MTH
    CLASS CORE ;
    FOREIGN NAND2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.825 1.540 1.965 ;
        RECT  1.250 0.825 1.330 0.985 ;
        RECT  0.935 1.805 1.330 1.965 ;
        RECT  0.990 0.385 1.250 0.985 ;
        RECT  0.675 1.805 0.935 2.405 ;
        END
        AntennaDiffArea 0.575 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.195 0.545 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 1.180 1.150 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.130 1.640 0.130 ;
        RECT  0.125 -0.130 0.385 1.010 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 2.740 1.640 3.000 ;
        RECT  1.215 2.145 1.475 3.000 ;
        RECT  0.385 2.740 1.215 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND2X2MTH

MACRO NAND2X3MTH
    CLASS CORE ;
    FOREIGN NAND2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 1.760 1.950 2.400 ;
        RECT  0.935 1.760 1.640 1.920 ;
        RECT  0.935 0.810 1.250 0.970 ;
        RECT  0.775 0.810 0.935 2.295 ;
        RECT  0.675 1.695 0.775 2.295 ;
        END
        AntennaDiffArea 0.68 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 0.905 2.080 1.425 ;
        RECT  1.590 0.905 1.820 1.065 ;
        RECT  1.430 0.470 1.590 1.065 ;
        RECT  0.595 0.470 1.430 0.630 ;
        RECT  0.435 0.470 0.595 1.480 ;
        RECT  0.100 0.880 0.435 1.480 ;
        END
        AntennaGateArea 0.286 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.115 1.245 1.540 1.580 ;
        END
        AntennaGateArea 0.286 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 -0.130 2.460 0.130 ;
        RECT  1.855 -0.130 2.115 0.725 ;
        RECT  0.385 -0.130 1.855 0.130 ;
        RECT  0.125 -0.130 0.385 0.295 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 2.460 3.000 ;
        RECT  0.125 1.740 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND2X3MTH

MACRO NAND2X4MTH
    CLASS CORE ;
    FOREIGN NAND2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 1.740 1.895 2.410 ;
        RECT  1.110 1.740 1.635 1.970 ;
        RECT  1.110 0.795 1.395 0.975 ;
        RECT  0.930 0.795 1.110 1.970 ;
        RECT  0.815 1.740 0.930 1.970 ;
        RECT  0.555 1.740 0.815 2.410 ;
        END
        AntennaDiffArea 0.98 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.935 0.880 1.985 1.510 ;
        RECT  1.825 0.455 1.935 1.510 ;
        RECT  1.775 0.455 1.825 1.040 ;
        RECT  0.750 0.455 1.775 0.615 ;
        RECT  0.590 0.455 0.750 1.540 ;
        RECT  0.310 1.205 0.590 1.540 ;
        RECT  0.100 1.205 0.310 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.155 1.635 1.560 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.330 -0.130 2.460 0.130 ;
        RECT  2.115 -0.130 2.330 0.700 ;
        RECT  0.410 -0.130 2.115 0.130 ;
        RECT  0.150 -0.130 0.410 1.025 ;
        RECT  0.000 -0.130 0.150 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.355 2.740 2.460 3.000 ;
        RECT  1.095 2.150 1.355 3.000 ;
        RECT  0.000 2.740 1.095 3.000 ;
        END
    END VDD
END NAND2X4MTH

MACRO NAND2X5MTH
    CLASS CORE ;
    FOREIGN NAND2X5MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.330 0.370 3.590 1.990 ;
        RECT  2.545 0.370 3.330 0.580 ;
        RECT  3.025 1.760 3.330 1.990 ;
        RECT  2.765 1.760 3.025 2.360 ;
        RECT  1.995 1.760 2.765 1.970 ;
        RECT  2.285 0.370 2.545 0.725 ;
        RECT  1.735 1.760 1.995 2.360 ;
        RECT  0.935 1.760 1.735 1.970 ;
        RECT  0.675 1.760 0.935 2.360 ;
        END
        AntennaDiffArea 1.276 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.615 1.275 1.555 1.540 ;
        END
        AntennaGateArea 0.5187 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.275 3.115 1.540 ;
        END
        AntennaGateArea 0.5187 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 -0.130 3.690 0.130 ;
        RECT  1.225 -0.130 1.485 0.675 ;
        RECT  0.385 -0.130 1.225 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 2.740 3.690 3.000 ;
        RECT  3.305 2.170 3.565 3.000 ;
        RECT  2.510 2.740 3.305 3.000 ;
        RECT  2.250 2.150 2.510 3.000 ;
        RECT  1.465 2.740 2.250 3.000 ;
        RECT  1.205 2.150 1.465 3.000 ;
        RECT  0.385 2.740 1.205 3.000 ;
        RECT  0.125 1.755 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.795 0.760 3.055 1.065 ;
        RECT  2.035 0.905 2.795 1.065 ;
        RECT  1.775 0.600 2.035 1.065 ;
        RECT  0.935 0.905 1.775 1.065 ;
        RECT  0.675 0.600 0.935 1.065 ;
    END
END NAND2X5MTH

MACRO NAND2X6MTH
    CLASS CORE ;
    FOREIGN NAND2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.290 0.345 3.560 2.030 ;
        RECT  2.250 0.345 3.290 0.615 ;
        RECT  3.025 1.700 3.290 2.030 ;
        RECT  2.970 1.700 3.025 2.370 ;
        RECT  2.765 1.760 2.970 2.370 ;
        RECT  1.995 1.760 2.765 2.030 ;
        RECT  1.735 1.760 1.995 2.375 ;
        RECT  0.935 1.760 1.735 2.030 ;
        RECT  0.675 1.760 0.935 2.380 ;
        END
        AntennaDiffArea 1.521 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.610 1.210 1.550 1.540 ;
        END
        AntennaGateArea 0.6162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 1.210 3.105 1.470 ;
        RECT  2.060 1.210 2.575 1.540 ;
        END
        AntennaGateArea 0.6162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.465 -0.130 3.690 0.130 ;
        RECT  1.205 -0.130 1.465 0.615 ;
        RECT  0.385 -0.130 1.205 0.130 ;
        RECT  0.125 -0.130 0.385 0.985 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 2.740 3.690 3.000 ;
        RECT  3.305 2.210 3.565 3.000 ;
        RECT  2.510 2.740 3.305 3.000 ;
        RECT  2.250 2.210 2.510 3.000 ;
        RECT  1.465 2.740 2.250 3.000 ;
        RECT  1.205 2.210 1.465 3.000 ;
        RECT  0.385 2.740 1.205 3.000 ;
        RECT  0.125 1.805 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.995 0.795 3.025 0.955 ;
        RECT  1.735 0.355 1.995 0.955 ;
        RECT  0.935 0.795 1.735 0.955 ;
        RECT  0.675 0.355 0.935 0.955 ;
    END
END NAND2X6MTH

MACRO NAND2X8MTH
    CLASS CORE ;
    FOREIGN NAND2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.120 0.470 4.410 1.925 ;
        RECT  1.185 0.470 4.120 0.770 ;
        RECT  3.880 1.575 4.120 1.925 ;
        RECT  3.530 1.575 3.880 2.490 ;
        RECT  2.955 1.905 3.530 2.255 ;
        RECT  2.575 1.905 2.955 2.505 ;
        RECT  1.985 1.905 2.575 2.255 ;
        RECT  1.605 1.865 1.985 2.465 ;
        RECT  0.960 1.865 1.605 2.125 ;
        RECT  0.580 1.865 0.960 2.465 ;
        END
        AntennaDiffArea 1.876 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.695 0.990 3.925 1.395 ;
        RECT  2.535 0.990 3.695 1.150 ;
        RECT  1.935 0.990 2.535 1.345 ;
        RECT  0.855 0.990 1.935 1.150 ;
        RECT  0.695 0.990 0.855 1.580 ;
        RECT  0.305 1.195 0.695 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.050 1.330 3.310 1.685 ;
        RECT  1.635 1.525 3.050 1.685 ;
        RECT  1.035 1.330 1.635 1.685 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  3.785 -0.130 4.385 0.290 ;
        RECT  2.325 -0.130 3.785 0.130 ;
        RECT  2.065 -0.130 2.325 0.290 ;
        RECT  0.515 -0.130 2.065 0.130 ;
        RECT  0.255 -0.130 0.515 0.980 ;
        RECT  0.000 -0.130 0.255 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 2.105 4.385 3.000 ;
        RECT  1.415 2.740 4.125 3.000 ;
        RECT  1.155 2.305 1.415 3.000 ;
        RECT  0.385 2.740 1.155 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND2X8MTH

MACRO NAND2XLMTH
    CLASS CORE ;
    FOREIGN NAND2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 0.765 1.540 1.920 ;
        RECT  1.135 0.765 1.325 1.025 ;
        RECT  0.685 1.760 1.325 1.920 ;
        END
        AntennaDiffArea 0.242 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.620 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.800 1.205 1.145 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.165 -0.130 1.640 0.130 ;
        RECT  0.485 -0.130 1.165 0.300 ;
        RECT  0.225 -0.130 0.485 1.025 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.490 2.740 1.640 3.000 ;
        RECT  1.230 2.100 1.490 3.000 ;
        RECT  0.945 2.740 1.230 3.000 ;
        RECT  0.685 2.570 0.945 3.000 ;
        RECT  0.385 2.740 0.685 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND2XLMTH

MACRO NAND3BX1MTH
    CLASS CORE ;
    FOREIGN NAND3BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.455 2.360 2.175 ;
        RECT  1.935 0.455 2.200 0.655 ;
        RECT  2.150 1.700 2.200 2.175 ;
        RECT  2.070 1.915 2.150 2.175 ;
        RECT  1.365 1.915 2.070 2.075 ;
        RECT  1.105 1.915 1.365 2.175 ;
        END
        AntennaDiffArea 0.575 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.195 1.150 1.735 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.290 1.915 1.680 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.390 1.545 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.015 -0.130 2.460 0.130 ;
        RECT  0.755 -0.130 1.015 0.335 ;
        RECT  0.000 -0.130 0.755 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.075 2.740 2.460 3.000 ;
        RECT  1.135 2.565 2.075 3.000 ;
        RECT  0.815 2.740 1.135 3.000 ;
        RECT  0.215 2.205 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.765 0.835 2.020 1.095 ;
        RECT  0.730 0.835 1.765 0.995 ;
        RECT  0.570 0.515 0.730 1.895 ;
        RECT  0.165 0.515 0.570 0.675 ;
        RECT  0.125 1.735 0.570 1.895 ;
    END
END NAND3BX1MTH

MACRO NAND3BX2MTH
    CLASS CORE ;
    FOREIGN NAND3BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.410 2.370 2.395 ;
        RECT  2.100 0.410 2.210 1.010 ;
        RECT  2.070 1.700 2.210 2.395 ;
        RECT  1.365 1.795 2.070 1.955 ;
        RECT  1.105 1.795 1.365 2.395 ;
        END
        AntennaDiffArea 0.92 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 0.880 1.150 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.880 1.580 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.380 1.625 ;
        END
        AntennaGateArea 0.0871 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 -0.130 2.460 0.130 ;
        RECT  0.310 -0.130 0.910 0.320 ;
        RECT  0.000 -0.130 0.310 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.805 2.740 2.460 3.000 ;
        RECT  0.205 2.315 0.805 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.920 1.225 2.030 1.485 ;
        RECT  1.760 0.540 1.920 1.485 ;
        RECT  0.720 0.540 1.760 0.700 ;
        RECT  0.560 0.540 0.720 1.965 ;
        RECT  0.125 0.815 0.560 0.975 ;
        RECT  0.125 1.805 0.560 1.965 ;
    END
END NAND3BX2MTH

MACRO NAND3BX4MTH
    CLASS CORE ;
    FOREIGN NAND3BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.785 4.000 2.395 ;
        RECT  2.475 0.785 3.790 0.965 ;
        RECT  3.520 2.215 3.790 2.395 ;
        RECT  3.260 2.215 3.520 2.475 ;
        RECT  2.430 2.215 3.260 2.395 ;
        RECT  2.260 0.365 2.475 0.965 ;
        RECT  2.170 2.215 2.430 2.475 ;
        RECT  1.475 2.215 2.170 2.395 ;
        RECT  1.215 2.215 1.475 2.475 ;
        END
        AntennaDiffArea 1.348 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 1.210 3.610 2.035 ;
        RECT  1.295 1.875 3.380 2.035 ;
        RECT  1.135 1.210 1.295 2.035 ;
        RECT  1.035 1.210 1.135 1.470 ;
        END
        AntennaGateArea 0.4108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.210 3.180 1.695 ;
        RECT  1.740 1.535 2.910 1.695 ;
        RECT  1.520 1.210 1.740 1.695 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.210 0.485 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.875 -0.130 4.100 0.130 ;
        RECT  3.615 -0.130 3.875 0.605 ;
        RECT  1.055 -0.130 3.615 0.130 ;
        RECT  0.795 -0.130 1.055 0.640 ;
        RECT  0.000 -0.130 0.795 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 2.740 4.100 3.000 ;
        RECT  2.710 2.575 2.970 3.000 ;
        RECT  0.925 2.740 2.710 3.000 ;
        RECT  0.665 2.110 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.080 1.195 2.645 1.355 ;
        RECT  1.920 0.820 2.080 1.355 ;
        RECT  0.825 0.820 1.920 0.980 ;
        RECT  0.665 0.820 0.825 1.920 ;
        RECT  0.515 0.820 0.665 0.980 ;
        RECT  0.385 1.760 0.665 1.920 ;
        RECT  0.255 0.610 0.515 0.980 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END NAND3BX4MTH

MACRO NAND3BXLMTH
    CLASS CORE ;
    FOREIGN NAND3BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.710 2.360 2.005 ;
        RECT  1.985 0.710 2.200 0.970 ;
        RECT  1.985 1.690 2.200 2.005 ;
        RECT  1.125 1.760 1.985 1.920 ;
        END
        AntennaDiffArea 0.367 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.195 1.300 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.110 2.110 1.655 2.360 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.100 0.400 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 -0.130 2.460 0.130 ;
        RECT  0.755 -0.130 1.695 0.355 ;
        RECT  0.000 -0.130 0.755 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.300 2.740 2.460 3.000 ;
        RECT  1.360 2.570 2.300 3.000 ;
        RECT  1.105 2.740 1.360 3.000 ;
        RECT  0.165 2.570 1.105 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.775 1.165 2.010 1.425 ;
        RECT  1.615 0.855 1.775 1.425 ;
        RECT  0.740 0.855 1.615 1.015 ;
        RECT  0.580 0.760 0.740 1.920 ;
        RECT  0.165 0.760 0.580 0.920 ;
        RECT  0.125 1.760 0.580 1.920 ;
    END
END NAND3BXLMTH

MACRO NAND3X12MTH
    CLASS CORE ;
    FOREIGN NAND3X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.255 1.720 9.665 2.390 ;
        RECT  7.485 0.785 9.645 1.110 ;
        RECT  8.615 1.720 9.255 2.125 ;
        RECT  8.175 1.720 8.615 2.380 ;
        RECT  7.540 1.720 8.175 2.125 ;
        RECT  7.485 1.720 7.540 2.380 ;
        RECT  7.040 0.785 7.485 2.380 ;
        RECT  6.865 0.785 7.040 2.125 ;
        RECT  6.035 1.720 6.865 2.125 ;
        RECT  4.570 1.720 6.035 2.400 ;
        RECT  3.905 1.720 4.570 2.125 ;
        RECT  2.570 1.720 3.905 2.400 ;
        RECT  1.935 1.720 2.570 2.125 ;
        RECT  0.585 1.720 1.935 2.415 ;
        END
        AntennaDiffArea 3.882 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.180 1.210 2.905 1.470 ;
        RECT  0.605 1.210 1.180 1.540 ;
        END
        AntennaGateArea 1.2324 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.490 1.210 6.050 1.470 ;
        RECT  4.045 1.210 4.490 1.540 ;
        RECT  3.410 1.210 4.045 1.470 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.560 1.330 9.775 1.490 ;
        RECT  7.815 1.330 8.560 1.540 ;
        END
        AntennaGateArea 1.2324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 -0.130 10.250 0.130 ;
        RECT  2.635 -0.130 2.895 0.565 ;
        RECT  0.905 -0.130 2.635 0.130 ;
        RECT  0.645 -0.130 0.905 0.570 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.115 2.740 10.250 3.000 ;
        RECT  9.855 1.865 10.115 3.000 ;
        RECT  9.065 2.740 9.855 3.000 ;
        RECT  8.805 2.315 9.065 3.000 ;
        RECT  7.990 2.740 8.805 3.000 ;
        RECT  7.730 2.305 7.990 3.000 ;
        RECT  6.845 2.740 7.730 3.000 ;
        RECT  6.245 2.355 6.845 3.000 ;
        RECT  4.365 2.740 6.245 3.000 ;
        RECT  4.105 2.305 4.365 3.000 ;
        RECT  2.375 2.740 4.105 3.000 ;
        RECT  2.115 2.305 2.375 3.000 ;
        RECT  0.385 2.740 2.115 3.000 ;
        RECT  0.125 1.830 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.855 0.405 10.115 0.975 ;
        RECT  3.675 0.405 9.855 0.565 ;
        RECT  3.425 0.750 6.485 0.910 ;
        RECT  3.165 0.410 3.425 0.910 ;
        RECT  2.375 0.750 3.165 0.910 ;
        RECT  2.115 0.410 2.375 0.910 ;
        RECT  1.425 0.750 2.115 0.910 ;
        RECT  1.165 0.410 1.425 0.910 ;
        RECT  0.390 0.750 1.165 0.910 ;
        RECT  0.130 0.410 0.390 0.910 ;
    END
END NAND3X12MTH

MACRO NAND3X1MTH
    CLASS CORE ;
    FOREIGN NAND3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.660 1.950 2.155 ;
        RECT  1.505 0.660 1.740 0.940 ;
        RECT  1.665 1.895 1.740 2.155 ;
        RECT  0.935 1.895 1.665 2.055 ;
        RECT  0.675 1.895 0.935 2.155 ;
        END
        AntennaDiffArea 0.577 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.160 0.635 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.815 1.145 1.130 1.715 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.120 1.560 1.715 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.705 -0.130 2.050 0.130 ;
        RECT  0.765 -0.130 1.705 0.300 ;
        RECT  0.425 -0.130 0.765 0.130 ;
        RECT  0.165 -0.130 0.425 0.980 ;
        RECT  0.000 -0.130 0.165 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.385 2.740 2.050 3.000 ;
        RECT  0.785 2.555 1.385 3.000 ;
        RECT  0.385 2.740 0.785 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3X1MTH

MACRO NAND3X2MTH
    CLASS CORE ;
    FOREIGN NAND3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.770 0.370 1.950 2.475 ;
        RECT  1.535 0.370 1.770 0.970 ;
        RECT  1.665 1.875 1.770 2.475 ;
        RECT  0.935 1.875 1.665 2.085 ;
        RECT  0.675 1.875 0.935 2.475 ;
        END
        AntennaDiffArea 0.881 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.645 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 0.880 1.130 1.575 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.150 1.575 1.695 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.435 -0.130 2.050 0.130 ;
        RECT  0.175 -0.130 0.435 0.980 ;
        RECT  0.000 -0.130 0.175 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 2.050 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3X2MTH

MACRO NAND3X3MTH
    CLASS CORE ;
    FOREIGN NAND3X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.515 3.590 1.710 ;
        RECT  1.765 0.515 3.380 0.675 ;
        RECT  3.125 1.550 3.380 1.710 ;
        RECT  2.965 1.550 3.125 2.220 ;
        RECT  0.675 2.060 2.965 2.220 ;
        END
        AntennaDiffArea 0.968 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 0.855 3.200 1.370 ;
        RECT  0.935 0.855 2.950 1.015 ;
        RECT  0.775 0.855 0.935 1.580 ;
        RECT  0.335 1.145 0.775 1.580 ;
        END
        AntennaGateArea 0.312 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.415 1.290 2.770 1.880 ;
        RECT  1.375 1.720 2.415 1.880 ;
        RECT  1.115 1.195 1.375 1.880 ;
        END
        AntennaGateArea 0.312 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 1.195 2.130 1.540 ;
        END
        AntennaGateArea 0.312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 -0.130 3.690 0.130 ;
        RECT  3.085 -0.130 3.345 0.335 ;
        RECT  0.595 -0.130 3.085 0.130 ;
        RECT  0.335 -0.130 0.595 0.865 ;
        RECT  0.000 -0.130 0.335 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 2.740 3.690 3.000 ;
        RECT  3.305 1.890 3.565 3.000 ;
        RECT  1.485 2.740 3.305 3.000 ;
        RECT  1.225 2.435 1.485 3.000 ;
        RECT  0.385 2.740 1.225 3.000 ;
        RECT  0.125 1.860 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3X3MTH

MACRO NAND3X4MTH
    CLASS CORE ;
    FOREIGN NAND3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.430 3.590 1.755 ;
        RECT  1.765 0.430 3.380 0.610 ;
        RECT  3.130 1.575 3.380 1.755 ;
        RECT  2.950 1.575 3.130 2.320 ;
        RECT  2.755 1.760 2.950 2.320 ;
        RECT  0.675 2.060 2.755 2.320 ;
        END
        AntennaDiffArea 1.412 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 0.790 3.200 1.395 ;
        RECT  0.835 0.790 3.040 0.950 ;
        RECT  0.675 0.790 0.835 1.580 ;
        RECT  0.335 1.160 0.675 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.575 1.210 2.770 1.580 ;
        RECT  2.415 1.210 2.575 1.880 ;
        RECT  1.275 1.720 2.415 1.880 ;
        RECT  1.015 1.205 1.275 1.880 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.595 1.205 2.195 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.460 -0.130 3.690 0.130 ;
        RECT  3.200 -0.130 3.460 0.250 ;
        RECT  0.495 -0.130 3.200 0.130 ;
        RECT  0.235 -0.130 0.495 0.980 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.570 2.740 3.690 3.000 ;
        RECT  3.310 1.935 3.570 3.000 ;
        RECT  1.485 2.740 3.310 3.000 ;
        RECT  1.225 2.505 1.485 3.000 ;
        RECT  0.385 2.740 1.225 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3X4MTH

MACRO NAND3X6MTH
    CLASS CORE ;
    FOREIGN NAND3X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 0.430 4.820 2.525 ;
        RECT  4.585 0.430 4.610 0.805 ;
        RECT  4.525 1.815 4.610 2.525 ;
        RECT  1.635 0.430 4.585 0.590 ;
        RECT  0.675 2.255 4.525 2.525 ;
        END
        AntennaDiffArea 2.133 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 0.770 3.255 1.395 ;
        RECT  0.855 0.770 3.095 0.930 ;
        RECT  0.695 0.770 0.855 1.580 ;
        RECT  0.395 1.160 0.695 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 1.315 3.950 2.075 ;
        RECT  2.545 1.915 3.790 2.075 ;
        RECT  2.285 1.450 2.545 2.075 ;
        RECT  2.110 1.740 2.285 2.075 ;
        RECT  1.195 1.915 2.110 2.075 ;
        RECT  1.035 1.230 1.195 2.075 ;
        END
        AntennaGateArea 0.6045 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.270 0.975 4.430 1.485 ;
        RECT  3.595 0.975 4.270 1.135 ;
        RECT  3.435 0.975 3.595 1.735 ;
        RECT  2.915 1.575 3.435 1.735 ;
        RECT  2.755 1.110 2.915 1.735 ;
        RECT  2.015 1.110 2.755 1.270 ;
        RECT  1.465 1.110 2.015 1.580 ;
        END
        AntennaGateArea 0.6045 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 -0.130 4.920 0.130 ;
        RECT  3.040 -0.130 3.300 0.250 ;
        RECT  0.505 -0.130 3.040 0.130 ;
        RECT  0.345 -0.130 0.505 0.980 ;
        RECT  0.000 -0.130 0.345 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 4.920 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3X6MTH

MACRO NAND3X8MTH
    CLASS CORE ;
    FOREIGN NAND3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.980 0.435 6.330 1.840 ;
        RECT  2.000 0.435 5.980 0.715 ;
        RECT  5.875 1.490 5.980 1.840 ;
        RECT  5.430 1.490 5.875 2.495 ;
        RECT  0.935 2.130 5.430 2.420 ;
        RECT  0.675 1.910 0.935 2.510 ;
        END
        AntennaDiffArea 1.958 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.640 0.895 5.800 1.225 ;
        RECT  3.605 0.895 5.640 1.055 ;
        RECT  3.005 0.895 3.605 1.270 ;
        RECT  0.755 0.895 3.005 1.055 ;
        RECT  0.370 0.895 0.755 1.605 ;
        END
        AntennaGateArea 0.624 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.080 1.235 5.270 1.395 ;
        RECT  3.920 1.235 4.080 1.610 ;
        RECT  2.770 1.450 3.920 1.610 ;
        RECT  2.490 1.235 2.770 1.610 ;
        RECT  1.610 1.235 2.490 1.395 ;
        RECT  1.350 1.235 1.610 1.465 ;
        END
        AntennaGateArea 0.624 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.480 1.575 4.860 1.950 ;
        RECT  2.090 1.790 4.480 1.950 ;
        RECT  1.830 1.575 2.090 1.950 ;
        END
        AntennaGateArea 0.624 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.060 -0.130 6.560 0.130 ;
        RECT  5.800 -0.130 6.060 0.250 ;
        RECT  3.440 -0.130 5.800 0.130 ;
        RECT  3.180 -0.130 3.440 0.250 ;
        RECT  0.935 -0.130 3.180 0.130 ;
        RECT  0.675 -0.130 0.935 0.715 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.425 2.740 6.560 3.000 ;
        RECT  6.165 2.045 6.425 3.000 ;
        RECT  2.430 2.740 6.165 3.000 ;
        RECT  2.170 2.620 2.430 3.000 ;
        RECT  0.385 2.740 2.170 3.000 ;
        RECT  0.125 2.050 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3X8MTH

MACRO NAND3XLMTH
    CLASS CORE ;
    FOREIGN NAND3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.705 1.950 1.930 ;
        RECT  1.545 0.705 1.740 0.965 ;
        RECT  0.675 1.770 1.740 1.930 ;
        END
        AntennaDiffArea 0.384 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.160 0.795 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.620 2.110 1.130 2.400 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 1.145 1.560 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.850 -0.130 2.050 0.130 ;
        RECT  0.910 -0.130 1.850 0.300 ;
        RECT  0.575 -0.130 0.910 0.130 ;
        RECT  0.315 -0.130 0.575 0.980 ;
        RECT  0.000 -0.130 0.315 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.850 2.740 2.050 3.000 ;
        RECT  1.310 2.375 1.850 3.000 ;
        RECT  0.935 2.740 1.310 3.000 ;
        RECT  0.675 2.615 0.935 3.000 ;
        RECT  0.385 2.740 0.675 3.000 ;
        RECT  0.125 1.760 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND3XLMTH

MACRO NAND4BBX1MTH
    CLASS CORE ;
    FOREIGN NAND4BBX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 0.480 3.600 2.465 ;
        RECT  2.755 0.480 3.440 0.640 ;
        RECT  2.905 2.305 3.440 2.465 ;
        RECT  2.745 2.150 2.905 2.465 ;
        RECT  2.495 0.375 2.755 0.640 ;
        RECT  2.325 2.150 2.745 2.360 ;
        RECT  2.065 2.015 2.325 2.360 ;
        RECT  1.365 2.200 2.065 2.360 ;
        RECT  1.105 2.015 1.365 2.360 ;
        END
        AntennaDiffArea 0.592 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.280 1.235 1.765 ;
        END
        AntennaGateArea 0.1274 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.210 0.330 1.580 0.720 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 1.095 3.260 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.240 0.400 1.685 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.375 -0.130 3.690 0.130 ;
        RECT  3.115 -0.130 3.375 0.300 ;
        RECT  0.920 -0.130 3.115 0.130 ;
        RECT  0.320 -0.130 0.920 0.360 ;
        RECT  0.000 -0.130 0.320 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.815 2.740 3.690 3.000 ;
        RECT  0.555 2.345 0.815 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.085 1.760 3.245 2.125 ;
        RECT  2.705 1.760 3.085 1.920 ;
        RECT  2.705 0.900 2.755 1.160 ;
        RECT  2.545 0.900 2.705 1.920 ;
        RECT  1.930 1.610 2.545 1.770 ;
        RECT  2.205 0.900 2.365 1.430 ;
        RECT  0.740 0.900 2.205 1.060 ;
        RECT  1.770 1.240 1.930 1.770 ;
        RECT  1.670 1.240 1.770 1.400 ;
        RECT  0.580 0.900 0.740 2.025 ;
        RECT  0.385 0.900 0.580 1.060 ;
        RECT  0.385 1.865 0.580 2.025 ;
        RECT  0.125 0.765 0.385 1.060 ;
        RECT  0.125 1.865 0.385 2.125 ;
    END
END NAND4BBX1MTH

MACRO NAND4BBX2MTH
    CLASS CORE ;
    FOREIGN NAND4BBX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.840 0.475 4.000 2.235 ;
        RECT  2.890 0.475 3.840 0.635 ;
        RECT  3.790 1.700 3.840 2.235 ;
        RECT  2.465 2.075 3.790 2.235 ;
        RECT  2.630 0.360 2.890 0.635 ;
        RECT  2.205 2.075 2.465 2.335 ;
        RECT  1.365 2.075 2.205 2.235 ;
        RECT  1.105 1.800 1.365 2.400 ;
        END
        AntennaDiffArea 0.99 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.150 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.955 1.565 1.605 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.300 1.155 3.660 1.540 ;
        END
        AntennaGateArea 0.0871 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.400 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.940 -0.130 4.100 0.130 ;
        RECT  3.340 -0.130 3.940 0.295 ;
        RECT  0.925 -0.130 3.340 0.130 ;
        RECT  0.325 -0.130 0.925 0.360 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.685 2.740 4.100 3.000 ;
        RECT  2.745 2.415 3.685 3.000 ;
        RECT  1.915 2.740 2.745 3.000 ;
        RECT  1.655 2.415 1.915 3.000 ;
        RECT  0.815 2.740 1.655 3.000 ;
        RECT  0.215 2.315 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.120 1.735 3.545 1.895 ;
        RECT  3.120 0.815 3.400 0.975 ;
        RECT  2.960 0.815 3.120 1.895 ;
        RECT  2.070 1.735 2.960 1.895 ;
        RECT  2.450 1.225 2.625 1.485 ;
        RECT  2.290 0.540 2.450 1.485 ;
        RECT  0.740 0.540 2.290 0.700 ;
        RECT  1.910 1.225 2.070 1.895 ;
        RECT  0.580 0.540 0.740 1.920 ;
        RECT  0.125 0.815 0.580 0.975 ;
        RECT  0.125 1.760 0.580 1.920 ;
    END
END NAND4BBX2MTH

MACRO NAND4BBX4MTH
    CLASS CORE ;
    FOREIGN NAND4BBX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.220 0.715 5.400 0.975 ;
        RECT  5.220 1.685 5.365 2.360 ;
        RECT  5.040 0.715 5.220 2.360 ;
        RECT  5.020 1.685 5.040 2.360 ;
        RECT  4.270 1.685 5.020 1.865 ;
        RECT  4.010 1.685 4.270 2.370 ;
        RECT  2.820 2.060 4.010 2.240 ;
        RECT  2.560 2.060 2.820 2.320 ;
        RECT  1.720 2.060 2.560 2.240 ;
        RECT  1.460 2.060 1.720 2.320 ;
        END
        AntennaDiffArea 1.612 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.260 1.990 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.380 1.260 2.980 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.090 1.105 0.380 1.600 ;
        END
        AntennaGateArea 0.1755 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.995 1.210 6.500 1.605 ;
        END
        AntennaGateArea 0.1755 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.335 -0.130 6.970 0.130 ;
        RECT  6.075 -0.130 6.335 0.615 ;
        RECT  0.380 -0.130 6.075 0.130 ;
        RECT  0.120 -0.130 0.380 0.925 ;
        RECT  0.000 -0.130 0.120 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.905 2.740 6.970 3.000 ;
        RECT  5.645 2.125 5.905 3.000 ;
        RECT  4.820 2.740 5.645 3.000 ;
        RECT  4.560 2.110 4.820 3.000 ;
        RECT  3.715 2.740 4.560 3.000 ;
        RECT  3.115 2.420 3.715 3.000 ;
        RECT  2.270 2.740 3.115 3.000 ;
        RECT  2.010 2.420 2.270 3.000 ;
        RECT  1.170 2.740 2.010 3.000 ;
        RECT  0.910 2.060 1.170 3.000 ;
        RECT  0.000 2.740 0.910 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.685 0.615 6.845 1.945 ;
        RECT  6.585 0.615 6.685 0.875 ;
        RECT  6.445 1.785 6.685 1.945 ;
        RECT  6.185 1.785 6.445 2.385 ;
        RECT  5.705 1.785 6.185 1.945 ;
        RECT  5.810 0.880 5.910 1.040 ;
        RECT  5.650 0.375 5.810 1.040 ;
        RECT  5.545 1.245 5.705 1.945 ;
        RECT  4.840 0.375 5.650 0.535 ;
        RECT  5.400 1.245 5.545 1.505 ;
        RECT  4.680 0.375 4.840 0.975 ;
        RECT  3.870 0.815 4.680 0.975 ;
        RECT  3.765 1.275 4.480 1.435 ;
        RECT  4.120 0.375 4.380 0.635 ;
        RECT  2.840 0.375 4.120 0.535 ;
        RECT  3.610 0.715 3.870 0.975 ;
        RECT  3.605 1.275 3.765 1.880 ;
        RECT  0.720 1.720 3.605 1.880 ;
        RECT  3.100 0.715 3.360 0.975 ;
        RECT  2.320 0.815 3.100 0.975 ;
        RECT  2.580 0.375 2.840 0.635 ;
        RECT  2.060 0.375 2.320 0.975 ;
        RECT  1.390 0.815 2.060 0.975 ;
        RECT  1.130 0.345 1.390 0.975 ;
        RECT  0.720 0.765 0.895 1.025 ;
        RECT  0.560 0.765 0.720 2.380 ;
        RECT  0.365 1.780 0.560 2.380 ;
    END
END NAND4BBX4MTH

MACRO NAND4BBXLMTH
    CLASS CORE ;
    FOREIGN NAND4BBXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.440 0.475 3.600 2.555 ;
        RECT  2.795 0.475 3.440 0.635 ;
        RECT  2.905 2.395 3.440 2.555 ;
        RECT  2.745 2.150 2.905 2.555 ;
        RECT  2.535 0.375 2.795 0.635 ;
        RECT  2.325 2.150 2.745 2.360 ;
        RECT  2.065 1.955 2.325 2.360 ;
        RECT  1.365 2.200 2.065 2.360 ;
        RECT  1.105 1.955 1.365 2.360 ;
        END
        AntennaDiffArea 0.382 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.290 1.235 1.765 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 0.330 1.660 0.720 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 1.095 3.260 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.390 1.775 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.375 -0.130 3.690 0.130 ;
        RECT  3.115 -0.130 3.375 0.290 ;
        RECT  0.925 -0.130 3.115 0.130 ;
        RECT  0.325 -0.130 0.925 0.360 ;
        RECT  0.000 -0.130 0.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 2.740 3.690 3.000 ;
        RECT  1.955 2.565 2.555 3.000 ;
        RECT  1.635 2.740 1.955 3.000 ;
        RECT  0.695 2.565 1.635 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.085 1.760 3.245 2.215 ;
        RECT  2.755 1.760 3.085 1.920 ;
        RECT  2.595 0.900 2.755 1.920 ;
        RECT  1.935 1.615 2.595 1.775 ;
        RECT  2.205 0.950 2.365 1.435 ;
        RECT  0.740 0.950 2.205 1.110 ;
        RECT  1.775 1.320 1.935 1.775 ;
        RECT  1.675 1.320 1.775 1.480 ;
        RECT  0.580 0.950 0.740 2.115 ;
        RECT  0.385 0.950 0.580 1.110 ;
        RECT  0.385 1.955 0.580 2.115 ;
        RECT  0.125 0.765 0.385 1.110 ;
        RECT  0.125 1.955 0.385 2.215 ;
    END
END NAND4BBXLMTH

MACRO NAND4BX1MTH
    CLASS CORE ;
    FOREIGN NAND4BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.480 2.770 2.030 ;
        RECT  2.475 0.480 2.610 0.740 ;
        RECT  2.560 1.700 2.610 2.030 ;
        RECT  2.330 1.870 2.560 2.030 ;
        RECT  2.070 1.870 2.330 2.130 ;
        RECT  1.365 1.870 2.070 2.030 ;
        RECT  1.105 1.870 1.365 2.130 ;
        END
        AntennaDiffArea 0.615 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.865 1.140 1.480 ;
        END
        AntennaGateArea 0.1274 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 1.030 1.540 1.655 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.720 0.865 1.955 1.495 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.400 1.500 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.975 -0.130 2.870 0.130 ;
        RECT  0.715 -0.130 0.975 0.345 ;
        RECT  0.000 -0.130 0.715 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.675 2.740 2.870 3.000 ;
        RECT  1.735 2.570 2.675 3.000 ;
        RECT  0.815 2.740 1.735 3.000 ;
        RECT  0.555 2.190 0.815 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.295 1.085 2.430 1.345 ;
        RECT  2.135 0.525 2.295 1.345 ;
        RECT  0.740 0.525 2.135 0.685 ;
        RECT  0.580 0.525 0.740 1.860 ;
        RECT  0.145 0.525 0.580 0.685 ;
        RECT  0.385 1.700 0.580 1.860 ;
        RECT  0.125 1.700 0.385 1.960 ;
    END
END NAND4BX1MTH

MACRO NAND4BX2MTH
    CLASS CORE ;
    FOREIGN NAND4BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.385 3.180 2.030 ;
        RECT  2.755 0.385 2.970 0.985 ;
        RECT  2.615 1.830 2.970 2.030 ;
        RECT  2.355 1.830 2.615 2.430 ;
        RECT  1.515 1.830 2.355 2.030 ;
        RECT  1.255 1.830 1.515 2.430 ;
        END
        AntennaDiffArea 0.923 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.150 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.350 1.770 1.580 ;
        RECT  1.330 1.045 1.560 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 0.880 2.235 1.470 ;
        RECT  1.740 0.880 1.950 1.170 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.165 0.400 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.990 -0.130 3.280 0.130 ;
        RECT  0.390 -0.130 0.990 0.360 ;
        RECT  0.000 -0.130 0.390 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.895 2.210 3.155 3.000 ;
        RECT  2.065 2.740 2.895 3.000 ;
        RECT  1.805 2.210 2.065 3.000 ;
        RECT  0.950 2.740 1.805 3.000 ;
        RECT  0.690 2.110 0.950 3.000 ;
        RECT  0.000 2.740 0.690 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.575 1.210 2.785 1.470 ;
        RECT  2.415 0.540 2.575 1.470 ;
        RECT  0.740 0.540 2.415 0.700 ;
        RECT  0.580 0.540 0.740 1.930 ;
        RECT  0.190 0.815 0.580 0.975 ;
        RECT  0.125 1.770 0.580 1.930 ;
    END
END NAND4BX2MTH

MACRO NAND4BX4MTH
    CLASS CORE ;
    FOREIGN NAND4BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.415 1.760 4.575 2.405 ;
        RECT  4.415 0.760 4.565 1.020 ;
        RECT  4.235 0.760 4.415 2.405 ;
        RECT  3.475 1.760 4.235 1.940 ;
        RECT  3.215 1.760 3.475 2.405 ;
        RECT  2.770 1.760 3.215 1.990 ;
        RECT  2.560 1.700 2.770 1.990 ;
        RECT  2.045 1.760 2.560 1.990 ;
        RECT  1.785 1.760 2.045 2.405 ;
        RECT  0.945 1.760 1.785 1.940 ;
        RECT  0.685 1.760 0.945 2.405 ;
        END
        AntennaDiffArea 1.634 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.495 1.210 1.130 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.210 2.160 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.070 1.210 3.670 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.285 1.190 5.685 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.485 -0.130 6.150 0.130 ;
        RECT  5.225 -0.130 5.485 0.545 ;
        RECT  0.925 -0.130 5.225 0.130 ;
        RECT  0.665 -0.130 0.925 0.615 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.120 2.740 6.150 3.000 ;
        RECT  4.860 2.100 5.120 3.000 ;
        RECT  4.025 2.740 4.860 3.000 ;
        RECT  3.765 2.120 4.025 3.000 ;
        RECT  2.760 2.740 3.765 3.000 ;
        RECT  2.500 2.170 2.760 3.000 ;
        RECT  1.495 2.740 2.500 3.000 ;
        RECT  1.235 2.120 1.495 3.000 ;
        RECT  0.395 2.740 1.235 3.000 ;
        RECT  0.135 1.830 0.395 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.865 0.615 6.025 1.920 ;
        RECT  5.765 0.615 5.865 0.875 ;
        RECT  5.660 1.760 5.865 1.920 ;
        RECT  5.400 1.760 5.660 2.360 ;
        RECT  4.915 1.760 5.400 1.920 ;
        RECT  4.975 0.765 5.075 1.025 ;
        RECT  4.815 0.405 4.975 1.025 ;
        RECT  4.755 1.210 4.915 1.920 ;
        RECT  4.055 0.405 4.815 0.565 ;
        RECT  4.595 1.210 4.755 1.470 ;
        RECT  3.795 0.405 4.055 0.955 ;
        RECT  2.755 0.795 3.795 0.955 ;
        RECT  1.725 0.355 3.535 0.615 ;
        RECT  1.465 0.795 2.505 0.955 ;
        RECT  1.205 0.355 1.465 0.955 ;
        RECT  0.385 0.795 1.205 0.955 ;
        RECT  0.125 0.355 0.385 0.955 ;
    END
END NAND4BX4MTH

MACRO NAND4BXLMTH
    CLASS CORE ;
    FOREIGN NAND4BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.675 2.770 1.990 ;
        RECT  2.480 0.675 2.610 0.935 ;
        RECT  2.560 1.700 2.610 1.990 ;
        RECT  1.105 1.770 2.560 1.930 ;
        END
        AntennaDiffArea 0.384 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.085 1.220 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.175 2.110 1.565 2.440 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 0.970 1.955 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.400 1.500 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 -0.130 2.870 0.130 ;
        RECT  1.905 -0.130 2.505 0.355 ;
        RECT  1.655 -0.130 1.905 0.130 ;
        RECT  0.715 -0.130 1.655 0.355 ;
        RECT  0.000 -0.130 0.715 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 2.740 2.870 3.000 ;
        RECT  1.805 2.570 2.745 3.000 ;
        RECT  1.495 2.740 1.805 3.000 ;
        RECT  0.815 2.620 1.495 3.000 ;
        RECT  0.555 2.230 0.815 3.000 ;
        RECT  0.000 2.740 0.555 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.295 1.165 2.430 1.425 ;
        RECT  2.135 0.540 2.295 1.425 ;
        RECT  0.740 0.540 2.135 0.700 ;
        RECT  0.580 0.540 0.740 1.845 ;
        RECT  0.145 0.540 0.580 0.700 ;
        RECT  0.385 1.685 0.580 1.845 ;
        RECT  0.125 1.685 0.385 1.945 ;
    END
END NAND4BXLMTH

MACRO NAND4X12MTH
    CLASS CORE ;
    FOREIGN NAND4X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.605 0.790 13.225 2.340 ;
        RECT  10.595 0.790 12.605 1.110 ;
        RECT  0.675 1.800 12.605 2.340 ;
        END
        AntennaDiffArea 4.86 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.540 1.275 3.180 1.580 ;
        END
        AntennaGateArea 1.2324 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.825 1.275 6.465 1.580 ;
        END
        AntennaGateArea 1.2324 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.005 1.275 9.985 1.580 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.465 1.330 12.425 1.540 ;
        END
        AntennaGateArea 1.2324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.060 -0.130 13.530 0.130 ;
        RECT  2.800 -0.130 3.060 0.565 ;
        RECT  1.990 -0.130 2.800 0.130 ;
        RECT  1.730 -0.130 1.990 0.565 ;
        RECT  0.920 -0.130 1.730 0.130 ;
        RECT  0.660 -0.130 0.920 0.565 ;
        RECT  0.000 -0.130 0.660 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 2.520 13.405 3.000 ;
        RECT  12.325 2.740 13.145 3.000 ;
        RECT  12.065 2.520 12.325 3.000 ;
        RECT  11.245 2.740 12.065 3.000 ;
        RECT  10.985 2.520 11.245 3.000 ;
        RECT  10.165 2.740 10.985 3.000 ;
        RECT  9.905 2.520 10.165 3.000 ;
        RECT  9.065 2.740 9.905 3.000 ;
        RECT  8.805 2.520 9.065 3.000 ;
        RECT  7.965 2.740 8.805 3.000 ;
        RECT  7.705 2.520 7.965 3.000 ;
        RECT  5.885 2.740 7.705 3.000 ;
        RECT  5.625 2.520 5.885 3.000 ;
        RECT  4.785 2.740 5.625 3.000 ;
        RECT  4.525 2.520 4.785 3.000 ;
        RECT  3.685 2.740 4.525 3.000 ;
        RECT  3.425 2.520 3.685 3.000 ;
        RECT  2.585 2.740 3.425 3.000 ;
        RECT  2.325 2.520 2.585 3.000 ;
        RECT  1.485 2.740 2.325 3.000 ;
        RECT  1.225 2.520 1.485 3.000 ;
        RECT  0.385 2.740 1.225 3.000 ;
        RECT  0.125 1.805 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.345 0.405 13.405 0.565 ;
        RECT  10.085 0.405 10.345 1.005 ;
        RECT  9.305 0.845 10.085 1.005 ;
        RECT  9.565 0.355 9.825 0.615 ;
        RECT  8.785 0.355 9.565 0.515 ;
        RECT  9.045 0.745 9.305 1.005 ;
        RECT  8.265 0.845 9.045 1.005 ;
        RECT  8.525 0.355 8.785 0.615 ;
        RECT  7.745 0.355 8.525 0.515 ;
        RECT  8.005 0.745 8.265 1.005 ;
        RECT  7.225 0.845 8.005 1.005 ;
        RECT  7.485 0.355 7.745 0.615 ;
        RECT  6.195 0.355 7.485 0.515 ;
        RECT  6.965 0.745 7.225 1.005 ;
        RECT  6.455 0.745 6.715 1.005 ;
        RECT  5.675 0.845 6.455 1.005 ;
        RECT  5.935 0.355 6.195 0.615 ;
        RECT  5.155 0.355 5.935 0.515 ;
        RECT  5.415 0.740 5.675 1.005 ;
        RECT  4.635 0.845 5.415 1.005 ;
        RECT  4.895 0.355 5.155 0.615 ;
        RECT  4.115 0.355 4.895 0.515 ;
        RECT  4.375 0.745 4.635 1.005 ;
        RECT  3.595 0.845 4.375 1.005 ;
        RECT  3.855 0.355 4.115 0.615 ;
        RECT  3.335 0.385 3.595 1.005 ;
        RECT  2.525 0.845 3.335 1.005 ;
        RECT  2.265 0.375 2.525 1.005 ;
        RECT  1.455 0.845 2.265 1.005 ;
        RECT  1.195 0.355 1.455 1.005 ;
        RECT  0.385 0.845 1.195 1.005 ;
        RECT  0.125 0.385 0.385 1.005 ;
    END
END NAND4X12MTH

MACRO NAND4X1MTH
    CLASS CORE ;
    FOREIGN NAND4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.660 2.360 1.930 ;
        RECT  1.865 0.660 2.150 0.920 ;
        RECT  0.555 1.770 2.150 1.930 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 1.205 0.675 1.465 ;
        RECT  0.100 1.205 0.355 1.580 ;
        END
        AntennaGateArea 0.1235 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.735 2.150 0.995 2.555 ;
        RECT  0.470 2.150 0.735 2.360 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.090 1.480 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.660 1.100 1.970 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 -0.130 2.460 0.130 ;
        RECT  0.985 -0.130 1.925 0.300 ;
        RECT  0.465 -0.130 0.985 0.130 ;
        RECT  0.205 -0.130 0.465 0.980 ;
        RECT  0.000 -0.130 0.205 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  2.075 2.230 2.335 3.000 ;
        RECT  1.775 2.740 2.075 3.000 ;
        RECT  1.175 2.570 1.775 3.000 ;
        RECT  0.385 2.740 1.175 3.000 ;
        RECT  0.125 2.570 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND4X1MTH

MACRO NAND4X2MTH
    CLASS CORE ;
    FOREIGN NAND4X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 0.440 2.365 1.990 ;
        RECT  1.985 0.440 2.205 0.700 ;
        RECT  2.150 1.700 2.205 1.990 ;
        RECT  1.915 1.810 2.150 1.990 ;
        RECT  1.655 1.810 1.915 2.410 ;
        RECT  0.935 1.810 1.655 1.990 ;
        RECT  0.675 1.810 0.935 2.410 ;
        END
        AntennaDiffArea 0.929 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.315 0.400 1.575 ;
        RECT  0.100 0.880 0.310 1.575 ;
        END
        AntennaGateArea 0.2054 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.815 0.880 1.110 1.480 ;
        RECT  0.510 0.880 0.815 1.170 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 0.880 1.560 1.480 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.880 2.025 1.480 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.425 -0.130 2.460 0.130 ;
        RECT  0.165 -0.130 0.425 0.700 ;
        RECT  0.000 -0.130 0.165 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 2.460 3.000 ;
        RECT  0.125 1.810 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND4X2MTH

MACRO NAND4X4MTH
    CLASS CORE ;
    FOREIGN NAND4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.660 2.305 3.835 2.465 ;
        RECT  0.740 0.405 2.355 0.565 ;
        RECT  0.580 0.405 0.740 1.065 ;
        RECT  0.500 2.275 0.660 2.465 ;
        RECT  0.260 0.905 0.580 1.065 ;
        RECT  0.310 2.275 0.500 2.435 ;
        RECT  0.260 2.110 0.310 2.435 ;
        RECT  0.100 0.905 0.260 2.435 ;
        END
        AntennaDiffArea 1.604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.925 1.220 4.025 1.480 ;
        RECT  3.765 1.220 3.925 2.125 ;
        RECT  1.195 1.965 3.765 2.125 ;
        RECT  1.035 1.755 1.195 2.125 ;
        RECT  0.720 1.755 1.035 1.915 ;
        RECT  0.440 1.245 0.720 1.915 ;
        END
        AntennaGateArea 0.4108 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 0.370 3.520 1.530 ;
        RECT  2.705 0.370 3.360 0.530 ;
        RECT  3.335 1.270 3.360 1.530 ;
        RECT  2.545 0.370 2.705 0.905 ;
        RECT  1.230 0.745 2.545 0.905 ;
        RECT  0.920 0.745 1.230 1.575 ;
        END
        AntennaGateArea 0.4108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 1.425 3.045 1.585 ;
        RECT  2.785 1.425 2.945 1.785 ;
        RECT  1.950 1.625 2.785 1.785 ;
        RECT  1.490 1.245 1.950 1.785 ;
        END
        AntennaGateArea 0.403 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.135 0.880 3.180 1.170 ;
        RECT  2.885 0.880 3.135 1.245 ;
        RECT  2.390 1.085 2.885 1.245 ;
        RECT  2.130 1.085 2.390 1.430 ;
        END
        AntennaGateArea 0.403 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.235 -0.130 4.510 0.130 ;
        RECT  3.975 -0.130 4.235 0.700 ;
        RECT  0.400 -0.130 3.975 0.130 ;
        RECT  0.240 -0.130 0.400 0.725 ;
        RECT  0.000 -0.130 0.240 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 1.890 4.385 3.000 ;
        RECT  0.385 2.740 4.125 3.000 ;
        RECT  0.125 2.615 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NAND4X4MTH

MACRO NAND4X6MTH
    CLASS CORE ;
    FOREIGN NAND4X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.450 0.345 6.720 2.075 ;
        RECT  5.440 0.345 6.450 0.615 ;
        RECT  6.300 1.290 6.450 2.075 ;
        RECT  6.250 1.290 6.300 2.405 ;
        RECT  6.040 1.805 6.250 2.405 ;
        RECT  5.275 1.805 6.040 2.075 ;
        RECT  5.015 1.805 5.275 2.405 ;
        RECT  4.175 1.805 5.015 2.075 ;
        RECT  3.915 1.805 4.175 2.405 ;
        RECT  3.075 1.805 3.915 2.075 ;
        RECT  2.815 1.805 3.075 2.405 ;
        RECT  1.975 1.805 2.815 2.075 ;
        RECT  1.715 1.805 1.975 2.405 ;
        RECT  0.935 1.805 1.715 2.075 ;
        RECT  0.675 1.805 0.935 2.405 ;
        END
        AntennaDiffArea 2.541 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.225 1.600 1.485 ;
        RECT  0.660 1.225 1.130 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 1.225 3.145 1.485 ;
        RECT  2.205 1.225 2.845 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.225 4.795 1.485 ;
        RECT  3.855 1.225 4.410 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.640 1.225 5.870 1.485 ;
        RECT  5.270 1.225 5.640 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.520 -0.130 6.970 0.130 ;
        RECT  1.260 -0.130 1.520 0.645 ;
        RECT  0.420 -0.130 1.260 0.130 ;
        RECT  0.160 -0.130 0.420 1.025 ;
        RECT  0.000 -0.130 0.160 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.840 2.740 6.970 3.000 ;
        RECT  6.580 2.255 6.840 3.000 ;
        RECT  5.790 2.740 6.580 3.000 ;
        RECT  5.530 2.255 5.790 3.000 ;
        RECT  4.725 2.740 5.530 3.000 ;
        RECT  4.465 2.255 4.725 3.000 ;
        RECT  3.625 2.740 4.465 3.000 ;
        RECT  3.365 2.255 3.625 3.000 ;
        RECT  2.525 2.740 3.365 3.000 ;
        RECT  2.265 2.255 2.525 3.000 ;
        RECT  1.455 2.740 2.265 3.000 ;
        RECT  1.195 2.255 1.455 3.000 ;
        RECT  0.385 2.740 1.195 3.000 ;
        RECT  0.125 1.805 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.950 0.795 6.210 0.985 ;
        RECT  5.190 0.825 5.950 0.985 ;
        RECT  4.930 0.385 5.190 0.985 ;
        RECT  4.150 0.825 4.930 0.985 ;
        RECT  4.410 0.385 4.670 0.645 ;
        RECT  3.630 0.385 4.410 0.545 ;
        RECT  3.890 0.725 4.150 0.985 ;
        RECT  3.370 0.385 3.630 0.985 ;
        RECT  2.590 0.385 3.370 0.545 ;
        RECT  2.850 0.725 3.110 0.985 ;
        RECT  2.070 0.825 2.850 0.985 ;
        RECT  2.330 0.385 2.590 0.645 ;
        RECT  1.810 0.385 2.070 0.985 ;
        RECT  0.970 0.825 1.810 0.985 ;
        RECT  0.710 0.385 0.970 0.985 ;
    END
END NAND4X6MTH

MACRO NAND4X8MTH
    CLASS CORE ;
    FOREIGN NAND4X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.765 0.785 8.795 1.125 ;
        RECT  8.505 0.785 8.765 2.400 ;
        RECT  8.300 0.785 8.505 2.150 ;
        RECT  7.515 0.785 8.300 1.125 ;
        RECT  7.685 1.800 8.300 2.150 ;
        RECT  7.425 1.800 7.685 2.400 ;
        RECT  6.595 1.800 7.425 2.150 ;
        RECT  6.335 1.800 6.595 2.400 ;
        RECT  5.495 1.800 6.335 2.150 ;
        RECT  5.235 1.800 5.495 2.400 ;
        RECT  4.235 1.800 5.235 2.150 ;
        RECT  3.975 1.800 4.235 2.400 ;
        RECT  3.135 1.800 3.975 2.150 ;
        RECT  2.875 1.800 3.135 2.400 ;
        RECT  2.035 1.800 2.875 2.150 ;
        RECT  1.775 1.800 2.035 2.400 ;
        RECT  0.935 1.800 1.775 2.150 ;
        RECT  0.675 1.800 0.935 2.400 ;
        END
        AntennaDiffArea 3.24 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.275 2.170 1.435 ;
        RECT  0.550 1.275 1.130 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.210 1.275 4.365 1.435 ;
        RECT  2.745 1.275 3.210 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.050 1.275 6.805 1.435 ;
        RECT  5.185 1.275 6.050 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.145 1.330 8.085 1.540 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 -0.130 9.430 0.130 ;
        RECT  1.785 -0.130 2.045 0.665 ;
        RECT  0.940 -0.130 1.785 0.130 ;
        RECT  0.680 -0.130 0.940 0.665 ;
        RECT  0.000 -0.130 0.680 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 2.740 9.430 3.000 ;
        RECT  9.045 1.800 9.305 3.000 ;
        RECT  8.225 2.740 9.045 3.000 ;
        RECT  7.965 2.330 8.225 3.000 ;
        RECT  7.145 2.740 7.965 3.000 ;
        RECT  6.885 2.330 7.145 3.000 ;
        RECT  6.045 2.740 6.885 3.000 ;
        RECT  5.785 2.330 6.045 3.000 ;
        RECT  4.865 2.740 5.785 3.000 ;
        RECT  4.605 2.330 4.865 3.000 ;
        RECT  3.685 2.740 4.605 3.000 ;
        RECT  3.425 2.330 3.685 3.000 ;
        RECT  2.585 2.740 3.425 3.000 ;
        RECT  2.325 2.330 2.585 3.000 ;
        RECT  1.485 2.740 2.325 3.000 ;
        RECT  1.225 2.330 1.485 3.000 ;
        RECT  0.385 2.740 1.225 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.045 0.405 9.305 1.005 ;
        RECT  7.265 0.405 9.045 0.565 ;
        RECT  7.005 0.375 7.265 1.005 ;
        RECT  6.225 0.845 7.005 1.005 ;
        RECT  6.485 0.385 6.745 0.645 ;
        RECT  5.705 0.385 6.485 0.545 ;
        RECT  5.965 0.745 6.225 1.005 ;
        RECT  5.185 0.845 5.965 1.005 ;
        RECT  5.445 0.385 5.705 0.645 ;
        RECT  4.155 0.385 5.445 0.545 ;
        RECT  4.925 0.745 5.185 1.005 ;
        RECT  4.415 0.745 4.675 1.005 ;
        RECT  3.635 0.845 4.415 1.005 ;
        RECT  3.895 0.385 4.155 0.645 ;
        RECT  3.115 0.385 3.895 0.545 ;
        RECT  3.375 0.745 3.635 1.005 ;
        RECT  2.595 0.845 3.375 1.005 ;
        RECT  2.855 0.385 3.115 0.645 ;
        RECT  2.335 0.385 2.595 1.005 ;
        RECT  1.495 0.845 2.335 1.005 ;
        RECT  1.235 0.385 1.495 1.005 ;
        RECT  0.385 0.845 1.235 1.005 ;
        RECT  0.125 0.385 0.385 1.005 ;
    END
END NAND4X8MTH

MACRO NAND4XLMTH
    CLASS CORE ;
    FOREIGN NAND4XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.720 2.360 1.920 ;
        RECT  1.945 0.720 2.150 0.980 ;
        RECT  0.585 1.760 2.150 1.920 ;
        END
        AntennaDiffArea 0.396 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 1.205 0.665 1.465 ;
        RECT  0.100 1.205 0.355 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 2.110 0.995 2.390 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.090 1.465 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.645 1.160 1.970 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 -0.130 2.460 0.130 ;
        RECT  1.530 -0.130 2.130 0.300 ;
        RECT  1.280 -0.130 1.530 0.130 ;
        RECT  0.680 -0.130 1.280 0.300 ;
        RECT  0.430 -0.130 0.680 0.130 ;
        RECT  0.170 -0.130 0.430 1.025 ;
        RECT  0.000 -0.130 0.170 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.250 2.740 2.460 3.000 ;
        RECT  1.310 2.570 2.250 3.000 ;
        RECT  1.130 2.740 1.310 3.000 ;
        RECT  0.190 2.570 1.130 3.000 ;
        RECT  0.000 2.740 0.190 3.000 ;
        END
    END VDD
END NAND4XLMTH

MACRO NOR2BX12MTH
    CLASS CORE ;
    FOREIGN NOR2BX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.770 0.435 8.070 2.440 ;
        RECT  7.265 0.435 7.770 1.375 ;
        RECT  2.735 1.935 7.770 2.440 ;
        RECT  2.205 0.435 7.265 0.805 ;
        END
        AntennaDiffArea 2.676 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.835 1.555 7.590 1.715 ;
        RECT  5.305 1.365 5.835 1.715 ;
        RECT  4.055 1.555 5.305 1.715 ;
        RECT  3.455 1.365 4.055 1.715 ;
        RECT  2.400 1.555 3.455 1.715 ;
        RECT  2.040 1.365 2.400 1.950 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.325 1.435 1.540 ;
        END
        AntennaGateArea 0.5304 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 -0.130 8.200 0.130 ;
        RECT  7.815 -0.130 8.075 0.250 ;
        RECT  5.020 -0.130 7.815 0.130 ;
        RECT  4.760 -0.130 5.020 0.250 ;
        RECT  1.945 -0.130 4.760 0.130 ;
        RECT  1.685 -0.130 1.945 0.795 ;
        RECT  0.925 -0.130 1.685 0.130 ;
        RECT  0.665 -0.130 0.925 0.795 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.700 2.740 8.200 3.000 ;
        RECT  7.100 2.620 7.700 3.000 ;
        RECT  5.620 2.740 7.100 3.000 ;
        RECT  5.360 2.620 5.620 3.000 ;
        RECT  3.870 2.740 5.360 3.000 ;
        RECT  3.610 2.620 3.870 3.000 ;
        RECT  2.115 2.740 3.610 3.000 ;
        RECT  1.855 2.130 2.115 3.000 ;
        RECT  1.035 2.740 1.855 3.000 ;
        RECT  0.775 2.140 1.035 3.000 ;
        RECT  0.000 2.740 0.775 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.305 1.025 6.670 1.345 ;
        RECT  4.880 1.025 6.305 1.185 ;
        RECT  4.395 1.025 4.880 1.345 ;
        RECT  3.180 1.025 4.395 1.185 ;
        RECT  2.580 1.025 3.180 1.345 ;
        RECT  1.850 1.025 2.580 1.185 ;
        RECT  1.690 0.985 1.850 1.880 ;
        RECT  1.435 0.985 1.690 1.145 ;
        RECT  1.575 1.720 1.690 1.880 ;
        RECT  1.315 1.720 1.575 2.360 ;
        RECT  1.175 0.660 1.435 1.145 ;
        RECT  0.495 1.720 1.315 1.880 ;
        RECT  0.415 0.985 1.175 1.145 ;
        RECT  0.235 1.720 0.495 2.335 ;
        RECT  0.155 0.660 0.415 1.145 ;
    END
END NOR2BX12MTH

MACRO NOR2BX1MTH
    CLASS CORE ;
    FOREIGN NOR2BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 0.920 1.950 2.125 ;
        RECT  1.470 0.920 1.790 1.080 ;
        RECT  1.650 1.700 1.790 2.125 ;
        RECT  1.310 0.540 1.470 1.080 ;
        RECT  1.155 0.540 1.310 0.800 ;
        END
        AntennaDiffArea 0.367 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.035 1.130 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.075 0.725 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 -0.130 2.050 0.130 ;
        RECT  1.665 -0.130 1.925 0.740 ;
        RECT  0.865 -0.130 1.665 0.130 ;
        RECT  0.265 -0.130 0.865 0.310 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 2.740 2.050 3.000 ;
        RECT  1.185 2.555 1.785 3.000 ;
        RECT  0.945 2.740 1.185 3.000 ;
        RECT  0.685 2.100 0.945 3.000 ;
        RECT  0.295 2.535 0.685 3.000 ;
        RECT  0.000 2.740 0.295 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.470 1.260 1.610 1.520 ;
        RECT  1.310 1.260 1.470 1.920 ;
        RECT  0.285 1.760 1.310 1.920 ;
        RECT  0.285 0.590 0.385 0.850 ;
        RECT  0.125 0.590 0.285 1.920 ;
    END
END NOR2BX1MTH

MACRO NOR2BX2MTH
    CLASS CORE ;
    FOREIGN NOR2BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 0.795 1.950 2.400 ;
        RECT  1.410 0.795 1.790 0.955 ;
        RECT  1.560 2.110 1.790 2.400 ;
        RECT  1.150 0.355 1.410 0.955 ;
        END
        AntennaDiffArea 0.57 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.135 1.260 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.450 1.155 0.740 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 -0.130 2.050 0.130 ;
        RECT  1.660 -0.130 1.920 0.615 ;
        RECT  0.855 -0.130 1.660 0.130 ;
        RECT  0.595 -0.130 0.855 0.460 ;
        RECT  0.000 -0.130 0.595 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 2.740 2.050 3.000 ;
        RECT  0.690 2.105 0.950 3.000 ;
        RECT  0.000 2.740 0.690 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.440 1.310 1.600 1.920 ;
        RECT  0.270 1.760 1.440 1.920 ;
        RECT  0.270 0.815 0.390 0.975 ;
        RECT  0.110 0.815 0.270 1.920 ;
    END
END NOR2BX2MTH

MACRO NOR2BX4MTH
    CLASS CORE ;
    FOREIGN NOR2BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.730 0.510 1.990 0.770 ;
        RECT  0.905 0.590 1.730 0.770 ;
        RECT  1.225 1.865 1.485 2.470 ;
        RECT  0.310 1.865 1.225 2.045 ;
        RECT  0.645 0.430 0.905 1.085 ;
        RECT  0.310 0.905 0.645 1.085 ;
        RECT  0.100 0.905 0.310 2.045 ;
        END
        AntennaDiffArea 0.968 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.310 2.115 1.685 ;
        RECT  0.785 1.525 1.955 1.685 ;
        RECT  0.490 1.275 0.785 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.295 1.290 2.770 1.605 ;
        END
        AntennaGateArea 0.1755 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.540 -0.130 3.280 0.130 ;
        RECT  2.280 -0.130 2.540 0.730 ;
        RECT  1.445 -0.130 2.280 0.130 ;
        RECT  1.185 -0.130 1.445 0.370 ;
        RECT  0.385 -0.130 1.185 0.130 ;
        RECT  0.125 -0.130 0.385 0.690 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.440 2.740 3.280 3.000 ;
        RECT  2.180 1.865 2.440 3.000 ;
        RECT  0.555 2.740 2.180 3.000 ;
        RECT  0.295 2.270 0.555 3.000 ;
        RECT  0.000 2.740 0.295 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.955 0.630 3.115 2.385 ;
        RECT  2.820 0.630 2.955 1.110 ;
        RECT  2.795 1.785 2.955 2.385 ;
        RECT  1.685 0.950 2.820 1.110 ;
        RECT  1.525 0.950 1.685 1.345 ;
        RECT  1.085 1.185 1.525 1.345 ;
    END
END NOR2BX4MTH

MACRO NOR2BX8MTH
    CLASS CORE ;
    FOREIGN NOR2BX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.015 0.430 3.965 0.730 ;
        RECT  3.045 1.905 3.395 2.505 ;
        RECT  1.490 1.905 3.045 2.255 ;
        RECT  0.905 0.350 3.015 0.730 ;
        RECT  1.140 1.905 1.490 2.505 ;
        RECT  0.380 1.905 1.140 2.255 ;
        RECT  0.585 0.350 0.905 1.095 ;
        RECT  0.380 0.745 0.585 1.095 ;
        RECT  0.100 0.745 0.380 2.255 ;
        END
        AntennaDiffArea 1.908 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 1.315 4.140 1.685 ;
        RECT  2.515 1.525 3.880 1.685 ;
        RECT  1.915 1.290 2.515 1.685 ;
        RECT  0.720 1.525 1.915 1.685 ;
        RECT  0.560 1.315 0.720 1.685 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.100 1.240 5.640 1.580 ;
        END
        AntennaGateArea 0.3536 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 1.025 ;
        RECT  4.525 -0.130 5.355 0.130 ;
        RECT  4.265 -0.130 4.525 0.740 ;
        RECT  3.425 -0.130 4.265 0.130 ;
        RECT  3.165 -0.130 3.425 0.250 ;
        RECT  0.390 -0.130 3.165 0.130 ;
        RECT  0.130 -0.130 0.390 0.565 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 2.740 5.740 3.000 ;
        RECT  5.355 1.795 5.615 3.000 ;
        RECT  4.565 2.740 5.355 3.000 ;
        RECT  3.965 1.865 4.565 3.000 ;
        RECT  2.325 2.740 3.965 3.000 ;
        RECT  2.065 2.440 2.325 3.000 ;
        RECT  0.525 2.740 2.065 3.000 ;
        RECT  0.265 2.480 0.525 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.915 1.760 5.105 2.360 ;
        RECT  4.915 0.580 5.075 0.840 ;
        RECT  4.755 0.580 4.915 2.360 ;
        RECT  3.480 0.950 4.755 1.110 ;
        RECT  2.880 0.950 3.480 1.345 ;
        RECT  1.570 0.950 2.880 1.110 ;
        RECT  1.410 0.950 1.570 1.345 ;
        RECT  1.205 1.185 1.410 1.345 ;
    END
END NOR2BX8MTH

MACRO NOR2BXLMTH
    CLASS CORE ;
    FOREIGN NOR2BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.790 0.735 1.950 2.030 ;
        RECT  1.175 0.735 1.790 0.895 ;
        RECT  1.670 1.690 1.790 2.030 ;
        END
        AntennaDiffArea 0.273 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 1.075 1.150 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.075 0.725 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.775 -0.130 2.050 0.130 ;
        RECT  0.835 -0.130 1.775 0.380 ;
        RECT  0.000 -0.130 0.835 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 2.740 2.050 3.000 ;
        RECT  1.240 2.620 1.840 3.000 ;
        RECT  0.970 2.740 1.240 3.000 ;
        RECT  0.710 2.100 0.970 3.000 ;
        RECT  0.000 2.740 0.710 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.490 1.170 1.610 1.430 ;
        RECT  1.330 1.170 1.490 1.920 ;
        RECT  0.285 1.760 1.330 1.920 ;
        RECT  0.285 0.735 0.385 0.895 ;
        RECT  0.125 0.735 0.285 1.920 ;
    END
END NOR2BXLMTH

MACRO NOR2X12MTH
    CLASS CORE ;
    FOREIGN NOR2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.930 0.500 6.370 2.440 ;
        RECT  5.635 0.500 5.930 1.375 ;
        RECT  4.710 2.000 5.930 2.440 ;
        RECT  4.955 0.500 5.635 1.000 ;
        RECT  4.580 0.355 4.955 1.000 ;
        RECT  4.450 1.935 4.710 2.440 ;
        RECT  1.620 0.355 4.580 0.805 ;
        RECT  2.990 2.000 4.450 2.440 ;
        RECT  2.730 1.935 2.990 2.440 ;
        RECT  1.270 2.000 2.730 2.440 ;
        RECT  0.645 0.355 1.620 0.740 ;
        RECT  1.010 1.935 1.270 2.440 ;
        END
        AntennaDiffArea 2.648 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.590 1.555 5.750 1.815 ;
        RECT  4.060 1.555 5.590 1.715 ;
        RECT  3.800 1.365 4.060 1.715 ;
        RECT  2.340 1.555 3.800 1.715 ;
        RECT  1.740 1.365 2.340 1.715 ;
        RECT  0.565 1.555 1.740 1.715 ;
        RECT  0.100 1.225 0.565 1.715 ;
        END
        AntennaGateArea 1.2324 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.400 1.185 4.815 1.345 ;
        RECT  4.240 1.025 4.400 1.345 ;
        RECT  3.135 1.025 4.240 1.185 ;
        RECT  2.875 1.025 3.135 1.345 ;
        RECT  1.440 1.025 2.875 1.185 ;
        RECT  0.840 0.920 1.440 1.345 ;
        END
        AntennaGateArea 1.2324 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.310 ;
        RECT  5.295 -0.130 6.175 0.130 ;
        RECT  5.135 -0.130 5.295 0.315 ;
        RECT  0.390 -0.130 5.135 0.130 ;
        RECT  0.130 -0.130 0.390 0.985 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.270 2.740 6.560 3.000 ;
        RECT  5.330 2.620 6.270 3.000 ;
        RECT  3.850 2.740 5.330 3.000 ;
        RECT  3.590 2.620 3.850 3.000 ;
        RECT  2.130 2.740 3.590 3.000 ;
        RECT  1.870 2.620 2.130 3.000 ;
        RECT  0.405 2.740 1.870 3.000 ;
        RECT  0.145 1.895 0.405 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
END NOR2X12MTH

MACRO NOR2X1MTH
    CLASS CORE ;
    FOREIGN NOR2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.765 1.275 2.360 ;
        RECT  0.755 0.715 0.915 2.360 ;
        END
        AntennaDiffArea 0.347 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.230 0.575 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.095 1.210 1.540 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 -0.130 1.640 0.130 ;
        RECT  1.245 -0.130 1.505 1.025 ;
        RECT  0.935 -0.130 1.245 0.130 ;
        RECT  0.675 -0.130 0.935 0.390 ;
        RECT  0.415 -0.130 0.675 0.130 ;
        RECT  0.155 -0.130 0.415 1.025 ;
        RECT  0.000 -0.130 0.155 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 2.740 1.640 3.000 ;
        RECT  0.415 2.620 1.105 3.000 ;
        RECT  0.155 1.765 0.415 3.000 ;
        RECT  0.000 2.740 0.155 3.000 ;
        END
    END VDD
END NOR2X1MTH

MACRO NOR2X2MTH
    CLASS CORE ;
    FOREIGN NOR2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.885 1.800 1.245 2.400 ;
        RECT  0.885 0.385 0.935 0.985 ;
        RECT  0.725 0.385 0.885 2.400 ;
        RECT  0.675 0.385 0.725 0.985 ;
        END
        AntennaDiffArea 0.57 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.515 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.065 1.225 1.540 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 -0.130 1.640 0.130 ;
        RECT  1.215 -0.130 1.475 1.025 ;
        RECT  0.385 -0.130 1.215 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 2.740 1.640 3.000 ;
        RECT  0.125 1.770 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NOR2X2MTH

MACRO NOR2X3MTH
    CLASS CORE ;
    FOREIGN NOR2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.580 2.360 2.025 ;
        RECT  2.150 0.580 2.200 1.170 ;
        RECT  1.400 1.865 2.200 2.025 ;
        RECT  0.795 0.580 2.150 0.740 ;
        RECT  1.140 1.865 1.400 2.125 ;
        RECT  0.535 0.580 0.795 0.890 ;
        END
        AntennaDiffArea 0.666 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.840 1.315 2.000 1.685 ;
        RECT  0.720 1.525 1.840 1.685 ;
        RECT  0.355 1.225 0.720 1.685 ;
        END
        AntennaGateArea 0.312 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.280 0.920 1.580 1.345 ;
        RECT  0.970 1.185 1.280 1.345 ;
        END
        AntennaGateArea 0.312 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.335 -0.130 2.460 0.130 ;
        RECT  1.075 -0.130 1.335 0.400 ;
        RECT  0.000 -0.130 1.075 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.260 2.740 2.460 3.000 ;
        RECT  2.000 2.210 2.260 3.000 ;
        RECT  0.540 2.740 2.000 3.000 ;
        RECT  0.280 1.875 0.540 3.000 ;
        RECT  0.000 2.740 0.280 3.000 ;
        END
    END VDD
END NOR2X3MTH

MACRO NOR2X4MTH
    CLASS CORE ;
    FOREIGN NOR2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.155 0.480 2.335 2.050 ;
        RECT  1.625 0.480 2.155 0.740 ;
        RECT  1.375 1.870 2.155 2.050 ;
        RECT  0.795 0.560 1.625 0.740 ;
        RECT  1.115 1.870 1.375 2.470 ;
        RECT  0.535 0.395 0.795 0.995 ;
        END
        AntennaDiffArea 0.878 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.815 1.225 1.975 1.685 ;
        RECT  0.720 1.525 1.815 1.685 ;
        RECT  0.355 1.225 0.720 1.685 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.170 0.920 1.580 1.345 ;
        RECT  0.945 1.185 1.170 1.345 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.340 -0.130 2.460 0.130 ;
        RECT  1.080 -0.130 1.340 0.380 ;
        RECT  0.000 -0.130 1.080 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 2.740 2.460 3.000 ;
        RECT  1.975 2.255 2.235 3.000 ;
        RECT  0.515 2.740 1.975 3.000 ;
        RECT  0.255 1.865 0.515 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
END NOR2X4MTH

MACRO NOR2X5MTH
    CLASS CORE ;
    FOREIGN NOR2X5MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.935 3.590 2.075 ;
        RECT  3.125 0.935 3.380 1.145 ;
        RECT  3.340 1.865 3.380 2.075 ;
        RECT  3.080 1.865 3.340 2.465 ;
        RECT  2.915 0.490 3.125 1.145 ;
        RECT  1.415 1.865 3.080 2.075 ;
        RECT  0.935 0.490 2.915 0.700 ;
        RECT  1.155 1.865 1.415 2.415 ;
        RECT  0.675 0.490 0.935 0.855 ;
        END
        AntennaDiffArea 1.282 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.260 2.385 1.685 ;
        RECT  0.735 1.525 1.740 1.685 ;
        RECT  0.475 1.225 0.735 1.685 ;
        END
        AntennaGateArea 0.5187 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.325 3.170 1.585 ;
        RECT  2.735 1.325 2.910 1.485 ;
        RECT  2.575 0.880 2.735 1.485 ;
        RECT  1.555 0.880 2.575 1.040 ;
        RECT  1.330 0.880 1.555 1.345 ;
        RECT  0.955 1.185 1.330 1.345 ;
        END
        AntennaGateArea 0.5187 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.675 ;
        RECT  2.480 -0.130 3.305 0.130 ;
        RECT  2.220 -0.130 2.480 0.300 ;
        RECT  0.385 -0.130 2.220 0.130 ;
        RECT  0.125 -0.130 0.385 1.000 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.385 2.740 3.690 3.000 ;
        RECT  2.125 2.325 2.385 3.000 ;
        RECT  0.525 2.740 2.125 3.000 ;
        RECT  0.265 1.915 0.525 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
END NOR2X5MTH

MACRO NOR2X6MTH
    CLASS CORE ;
    FOREIGN NOR2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.320 0.795 3.590 2.375 ;
        RECT  3.175 0.795 3.320 1.065 ;
        RECT  3.080 1.775 3.320 2.375 ;
        RECT  2.905 0.430 3.175 1.065 ;
        RECT  1.415 1.935 3.080 2.205 ;
        RECT  0.905 0.430 2.905 0.700 ;
        RECT  1.155 1.935 1.415 2.465 ;
        RECT  0.645 0.430 0.905 0.930 ;
        END
        AntennaDiffArea 1.52 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.260 2.385 1.735 ;
        RECT  0.685 1.575 1.740 1.735 ;
        RECT  0.525 1.225 0.685 1.735 ;
        END
        AntennaGateArea 0.6162 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 1.245 3.120 1.505 ;
        RECT  2.725 1.245 2.960 1.405 ;
        RECT  2.565 0.880 2.725 1.405 ;
        RECT  1.540 0.880 2.565 1.040 ;
        RECT  1.330 0.880 1.540 1.395 ;
        RECT  1.040 1.135 1.330 1.395 ;
        END
        AntennaGateArea 0.6162 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 -0.130 3.690 0.130 ;
        RECT  3.355 -0.130 3.515 0.615 ;
        RECT  2.480 -0.130 3.355 0.130 ;
        RECT  2.220 -0.130 2.480 0.250 ;
        RECT  0.390 -0.130 2.220 0.130 ;
        RECT  0.130 -0.130 0.390 0.985 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.385 2.740 3.690 3.000 ;
        RECT  2.125 2.385 2.385 3.000 ;
        RECT  0.525 2.740 2.125 3.000 ;
        RECT  0.265 1.915 0.525 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
END NOR2X6MTH

MACRO NOR2X8MTH
    CLASS CORE ;
    FOREIGN NOR2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.380 1.085 4.410 1.785 ;
        RECT  3.990 0.785 4.380 2.255 ;
        RECT  3.905 0.785 3.990 1.135 ;
        RECT  3.205 1.905 3.990 2.255 ;
        RECT  3.555 0.350 3.905 1.135 ;
        RECT  0.905 0.350 3.555 0.700 ;
        RECT  2.945 1.905 3.205 2.505 ;
        RECT  1.325 1.905 2.945 2.255 ;
        RECT  1.065 1.905 1.325 2.505 ;
        RECT  0.645 0.350 0.905 0.955 ;
        END
        AntennaDiffArea 1.756 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.645 1.315 3.805 1.685 ;
        RECT  2.405 1.525 3.645 1.685 ;
        RECT  1.760 1.290 2.405 1.685 ;
        RECT  0.625 1.525 1.760 1.685 ;
        RECT  0.465 1.225 0.625 1.685 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 1.185 3.375 1.345 ;
        RECT  2.665 0.920 2.825 1.345 ;
        RECT  1.580 0.920 2.665 1.080 ;
        RECT  1.285 0.920 1.580 1.345 ;
        RECT  0.895 1.185 1.285 1.345 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.345 -0.130 4.510 0.130 ;
        RECT  4.085 -0.130 4.345 0.605 ;
        RECT  0.390 -0.130 4.085 0.130 ;
        RECT  0.130 -0.130 0.390 0.985 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.215 2.740 4.510 3.000 ;
        RECT  3.955 2.570 4.215 3.000 ;
        RECT  2.205 2.740 3.955 3.000 ;
        RECT  1.945 2.570 2.205 3.000 ;
        RECT  0.465 2.740 1.945 3.000 ;
        RECT  0.205 1.915 0.465 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
END NOR2X8MTH

MACRO NOR2XLMTH
    CLASS CORE ;
    FOREIGN NOR2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.640 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.760 1.305 2.400 ;
        RECT  0.755 0.765 0.915 2.400 ;
        END
        AntennaDiffArea 0.238 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.230 0.575 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.095 1.210 1.540 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.505 -0.130 1.640 0.130 ;
        RECT  0.810 -0.130 1.505 0.510 ;
        RECT  0.385 -0.130 0.810 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 2.740 1.640 3.000 ;
        RECT  0.845 2.620 1.445 3.000 ;
        RECT  0.415 2.740 0.845 3.000 ;
        RECT  0.155 1.765 0.415 3.000 ;
        RECT  0.000 2.740 0.155 3.000 ;
        END
    END VDD
END NOR2XLMTH

MACRO NOR3BX1MTH
    CLASS CORE ;
    FOREIGN NOR3BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.755 2.360 2.175 ;
        RECT  1.105 0.755 2.200 0.915 ;
        RECT  2.065 1.700 2.200 2.175 ;
        END
        AntennaDiffArea 0.507 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.095 1.130 1.620 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.095 1.545 1.665 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.355 1.665 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.290 -0.130 2.460 0.130 ;
        RECT  2.030 -0.130 2.290 0.320 ;
        RECT  1.730 -0.130 2.030 0.130 ;
        RECT  0.790 -0.130 1.730 0.380 ;
        RECT  0.445 -0.130 0.790 0.130 ;
        RECT  0.185 -0.130 0.445 0.320 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.090 2.740 2.460 3.000 ;
        RECT  1.150 2.555 2.090 3.000 ;
        RECT  0.955 2.740 1.150 3.000 ;
        RECT  0.695 2.555 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.885 1.225 2.000 1.485 ;
        RECT  1.725 1.225 1.885 2.005 ;
        RECT  0.695 1.845 1.725 2.005 ;
        RECT  0.535 0.815 0.695 2.005 ;
        RECT  0.125 0.815 0.535 0.975 ;
        RECT  0.125 1.845 0.535 2.005 ;
    END
END NOR3BX1MTH

MACRO NOR3BX2MTH
    CLASS CORE ;
    FOREIGN NOR3BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.190 0.355 2.360 2.445 ;
        RECT  2.075 0.355 2.190 0.955 ;
        RECT  2.150 1.700 2.190 2.445 ;
        RECT  1.965 2.185 2.150 2.445 ;
        RECT  1.405 0.795 2.075 0.955 ;
        RECT  1.145 0.355 1.405 0.955 ;
        END
        AntennaDiffArea 0.807 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.885 1.135 1.130 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 1.135 1.630 1.660 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.355 1.665 ;
        END
        AntennaGateArea 0.0871 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 -0.130 2.460 0.130 ;
        RECT  0.265 -0.130 0.865 0.475 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.885 2.740 2.460 3.000 ;
        RECT  0.285 2.345 0.885 3.000 ;
        RECT  0.000 2.740 0.285 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.970 1.225 2.005 1.485 ;
        RECT  1.810 1.225 1.970 2.005 ;
        RECT  0.695 1.845 1.810 2.005 ;
        RECT  0.535 0.815 0.695 2.005 ;
        RECT  0.125 0.815 0.535 0.975 ;
        RECT  0.125 1.845 0.535 2.005 ;
    END
END NOR3BX2MTH

MACRO NOR3BX4MTH
    CLASS CORE ;
    FOREIGN NOR3BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.650 4.000 1.945 ;
        RECT  3.470 0.650 3.790 0.830 ;
        RECT  2.515 1.765 3.790 1.945 ;
        RECT  3.290 0.385 3.470 0.830 ;
        RECT  1.130 0.385 3.290 0.565 ;
        RECT  2.335 1.765 2.515 2.360 ;
        RECT  2.095 2.100 2.335 2.360 ;
        END
        AntennaDiffArea 1.216 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.305 1.025 3.565 1.445 ;
        RECT  3.110 1.025 3.305 1.185 ;
        RECT  2.950 0.745 3.110 1.185 ;
        RECT  1.275 0.745 2.950 0.905 ;
        RECT  1.115 0.745 1.275 1.515 ;
        RECT  0.920 0.875 1.115 1.515 ;
        END
        AntennaGateArea 0.403 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.365 3.085 1.580 ;
        RECT  2.560 1.085 2.770 1.580 ;
        RECT  1.615 1.085 2.560 1.245 ;
        RECT  1.455 1.085 1.615 1.455 ;
        END
        AntennaGateArea 0.403 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 0.985 0.720 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.100 0.130 ;
        RECT  3.715 -0.130 3.975 0.420 ;
        RECT  0.895 -0.130 3.715 0.130 ;
        RECT  0.635 -0.130 0.895 0.665 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.805 2.740 4.100 3.000 ;
        RECT  3.545 2.135 3.805 3.000 ;
        RECT  0.955 2.740 3.545 3.000 ;
        RECT  0.695 2.100 0.955 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.885 1.425 2.145 1.920 ;
        RECT  0.385 1.760 1.885 1.920 ;
        RECT  0.260 0.515 0.385 0.775 ;
        RECT  0.260 1.760 0.385 2.385 ;
        RECT  0.100 0.515 0.260 2.385 ;
    END
END NOR3BX4MTH

MACRO NOR3BXLMTH
    CLASS CORE ;
    FOREIGN NOR3BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.755 2.360 2.005 ;
        RECT  1.075 0.755 2.200 0.915 ;
        RECT  2.065 1.700 2.200 2.005 ;
        END
        AntennaDiffArea 0.399 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.095 1.130 1.620 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.095 1.545 1.665 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.040 0.355 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.230 -0.130 2.460 0.130 ;
        RECT  1.970 -0.130 2.230 0.300 ;
        RECT  1.660 -0.130 1.970 0.130 ;
        RECT  0.720 -0.130 1.660 0.380 ;
        RECT  0.000 -0.130 0.720 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 2.740 2.460 3.000 ;
        RECT  1.170 2.560 2.110 3.000 ;
        RECT  0.855 2.740 1.170 3.000 ;
        RECT  0.595 2.185 0.855 3.000 ;
        RECT  0.000 2.740 0.595 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.885 1.225 2.000 1.485 ;
        RECT  1.725 1.225 1.885 2.005 ;
        RECT  0.695 1.845 1.725 2.005 ;
        RECT  0.535 0.685 0.695 2.005 ;
        RECT  0.395 0.685 0.535 0.845 ;
        RECT  0.125 1.760 0.535 2.005 ;
        RECT  0.135 0.385 0.395 0.845 ;
    END
END NOR3BXLMTH

MACRO NOR3X12MTH
    CLASS CORE ;
    FOREIGN NOR3X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.505 1.495 9.125 2.440 ;
        RECT  6.040 0.310 8.785 0.565 ;
        RECT  7.305 1.865 8.505 2.440 ;
        RECT  5.235 2.205 7.305 2.440 ;
        RECT  4.525 0.310 6.040 0.590 ;
        RECT  4.180 1.905 5.235 2.440 ;
        RECT  3.905 0.430 4.525 0.590 ;
        RECT  1.885 2.205 4.180 2.440 ;
        RECT  3.360 0.310 3.905 0.590 ;
        RECT  1.045 0.310 3.360 0.565 ;
        RECT  0.325 2.060 1.885 2.440 ;
        RECT  0.605 0.310 1.045 0.905 ;
        RECT  0.325 0.530 0.605 0.905 ;
        RECT  0.090 0.530 0.325 2.440 ;
        END
        AntennaDiffArea 3.558 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.865 1.155 9.005 1.315 ;
        RECT  8.705 0.745 8.865 1.315 ;
        RECT  6.395 0.745 8.705 0.905 ;
        RECT  6.235 0.745 6.395 1.345 ;
        RECT  6.135 0.770 6.235 1.345 ;
        RECT  3.275 0.770 6.135 0.930 ;
        RECT  3.175 0.770 3.275 1.345 ;
        RECT  3.015 0.745 3.175 1.345 ;
        RECT  1.385 0.745 3.015 0.905 ;
        RECT  1.225 0.745 1.385 1.245 ;
        RECT  0.720 1.085 1.225 1.245 ;
        RECT  0.505 1.085 0.720 1.580 ;
        END
        AntennaGateArea 1.1895 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.045 1.155 8.525 1.315 ;
        RECT  7.885 1.155 8.045 1.685 ;
        RECT  7.225 1.525 7.885 1.685 ;
        RECT  7.125 1.425 7.225 1.685 ;
        RECT  6.965 1.425 7.125 2.025 ;
        RECT  5.615 1.865 6.965 2.025 ;
        RECT  5.455 1.450 5.615 2.025 ;
        RECT  5.355 1.450 5.455 1.685 ;
        RECT  4.085 1.525 5.355 1.685 ;
        RECT  3.955 1.450 4.085 1.685 ;
        RECT  3.825 1.450 3.955 2.025 ;
        RECT  3.795 1.490 3.825 2.025 ;
        RECT  2.495 1.865 3.795 2.025 ;
        RECT  2.235 1.425 2.495 2.025 ;
        RECT  2.110 1.720 2.235 2.025 ;
        RECT  1.195 1.720 2.110 1.880 ;
        RECT  0.935 1.425 1.195 1.880 ;
        END
        AntennaGateArea 1.1817 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.445 1.085 7.705 1.345 ;
        RECT  6.735 1.085 7.445 1.245 ;
        RECT  6.575 1.085 6.735 1.685 ;
        RECT  5.955 1.525 6.575 1.685 ;
        RECT  5.795 1.110 5.955 1.685 ;
        RECT  5.000 1.110 5.795 1.270 ;
        RECT  4.400 1.110 5.000 1.345 ;
        RECT  3.615 1.110 4.400 1.270 ;
        RECT  3.455 1.110 3.615 1.685 ;
        RECT  2.835 1.525 3.455 1.685 ;
        RECT  2.675 1.085 2.835 1.685 ;
        RECT  2.045 1.085 2.675 1.245 ;
        RECT  1.565 1.085 2.045 1.540 ;
        END
        AntennaGateArea 1.1817 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 -0.130 9.430 0.130 ;
        RECT  9.045 -0.130 9.305 0.955 ;
        RECT  4.345 -0.130 9.045 0.130 ;
        RECT  4.085 -0.130 4.345 0.250 ;
        RECT  0.385 -0.130 4.085 0.130 ;
        RECT  0.125 -0.130 0.385 0.305 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.215 2.740 9.430 3.000 ;
        RECT  8.955 2.620 9.215 3.000 ;
        RECT  6.505 2.740 8.955 3.000 ;
        RECT  6.245 2.620 6.505 3.000 ;
        RECT  3.215 2.740 6.245 3.000 ;
        RECT  2.955 2.620 3.215 3.000 ;
        RECT  0.500 2.740 2.955 3.000 ;
        RECT  0.240 2.620 0.500 3.000 ;
        RECT  0.000 2.740 0.240 3.000 ;
        END
    END VDD
END NOR3X12MTH

MACRO NOR3X1MTH
    CLASS CORE ;
    FOREIGN NOR3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.710 1.950 2.180 ;
        RECT  1.665 0.710 1.740 0.970 ;
        RECT  1.505 1.920 1.740 2.180 ;
        RECT  0.935 0.810 1.665 0.970 ;
        RECT  0.675 0.710 0.935 0.970 ;
        END
        AntennaDiffArea 0.473 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.585 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 1.155 1.130 1.825 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.155 1.550 1.740 ;
        END
        AntennaGateArea 0.1274 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.725 -0.130 2.050 0.130 ;
        RECT  0.785 -0.130 1.725 0.380 ;
        RECT  0.385 -0.130 0.785 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 2.740 2.050 3.000 ;
        RECT  0.715 2.570 1.655 3.000 ;
        RECT  0.425 2.740 0.715 3.000 ;
        RECT  0.165 1.770 0.425 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
END NOR3X1MTH

MACRO NOR3X2MTH
    CLASS CORE ;
    FOREIGN NOR3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.760 0.355 1.950 2.130 ;
        RECT  1.740 0.355 1.760 2.515 ;
        RECT  1.665 0.355 1.740 0.955 ;
        RECT  1.500 1.915 1.740 2.515 ;
        RECT  0.905 0.795 1.665 0.955 ;
        RECT  0.645 0.355 0.905 0.955 ;
        END
        AntennaDiffArea 0.813 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.625 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 1.180 1.130 1.905 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.170 1.560 1.705 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.390 -0.130 2.050 0.130 ;
        RECT  0.130 -0.130 0.390 0.955 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.445 2.740 2.050 3.000 ;
        RECT  0.185 1.785 0.445 3.000 ;
        RECT  0.000 2.740 0.185 3.000 ;
        END
    END VDD
END NOR3X2MTH

MACRO NOR3X4MTH
    CLASS CORE ;
    FOREIGN NOR3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.630 3.590 2.245 ;
        RECT  3.015 0.630 3.380 0.810 ;
        RECT  1.975 2.065 3.380 2.245 ;
        RECT  2.755 0.520 3.015 0.810 ;
        RECT  1.995 0.630 2.755 0.810 ;
        RECT  1.735 0.520 1.995 0.810 ;
        RECT  1.715 2.065 1.975 2.325 ;
        RECT  0.905 0.630 1.735 0.810 ;
        RECT  0.645 0.525 0.905 0.810 ;
        END
        AntennaDiffArea 1.288 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 0.990 3.185 1.485 ;
        RECT  0.735 0.990 2.925 1.150 ;
        RECT  0.575 0.990 0.735 1.580 ;
        RECT  0.405 1.225 0.575 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.445 1.365 2.705 1.885 ;
        RECT  1.250 1.725 2.445 1.885 ;
        RECT  0.920 1.365 1.250 1.990 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.545 1.330 2.180 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.565 -0.130 3.690 0.130 ;
        RECT  3.305 -0.130 3.565 0.450 ;
        RECT  1.455 -0.130 3.305 0.130 ;
        RECT  1.195 -0.130 1.455 0.450 ;
        RECT  0.390 -0.130 1.195 0.130 ;
        RECT  0.130 -0.130 0.390 0.955 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 2.740 3.690 3.000 ;
        RECT  3.135 2.430 3.395 3.000 ;
        RECT  0.590 2.740 3.135 3.000 ;
        RECT  0.330 1.915 0.590 3.000 ;
        RECT  0.000 2.740 0.330 3.000 ;
        END
    END VDD
END NOR3X4MTH

MACRO NOR3X6MTH
    CLASS CORE ;
    FOREIGN NOR3X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.585 0.405 4.830 2.440 ;
        RECT  4.535 0.405 4.585 0.905 ;
        RECT  4.175 1.765 4.585 2.440 ;
        RECT  3.805 0.745 4.535 0.905 ;
        RECT  1.815 2.260 4.175 2.440 ;
        RECT  3.435 0.310 3.805 0.905 ;
        RECT  0.645 0.310 3.435 0.565 ;
        RECT  1.555 2.160 1.815 2.440 ;
        END
        AntennaDiffArea 1.936 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.035 0.745 3.195 1.395 ;
        RECT  0.730 0.745 3.035 0.905 ;
        RECT  0.570 0.745 0.730 1.580 ;
        RECT  0.405 1.225 0.570 1.580 ;
        END
        AntennaGateArea 0.6006 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.875 1.425 3.975 1.585 ;
        RECT  3.715 1.425 3.875 2.080 ;
        RECT  2.465 1.920 3.715 2.080 ;
        RECT  2.205 1.425 2.465 2.080 ;
        RECT  1.165 1.720 2.205 1.880 ;
        RECT  0.920 1.315 1.165 1.990 ;
        END
        AntennaGateArea 0.6006 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 1.085 4.405 1.505 ;
        RECT  3.535 1.085 4.245 1.245 ;
        RECT  3.375 1.085 3.535 1.740 ;
        RECT  2.855 1.580 3.375 1.740 ;
        RECT  2.695 1.085 2.855 1.740 ;
        RECT  1.990 1.085 2.695 1.245 ;
        RECT  1.415 1.085 1.990 1.540 ;
        END
        AntennaGateArea 0.6006 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.285 -0.130 4.920 0.130 ;
        RECT  4.025 -0.130 4.285 0.565 ;
        RECT  0.390 -0.130 4.025 0.130 ;
        RECT  0.130 -0.130 0.390 0.955 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.185 2.740 4.920 3.000 ;
        RECT  2.925 2.620 3.185 3.000 ;
        RECT  0.510 2.740 2.925 3.000 ;
        RECT  0.250 1.915 0.510 3.000 ;
        RECT  0.000 2.740 0.250 3.000 ;
        END
    END VDD
END NOR3X6MTH

MACRO NOR3X8MTH
    CLASS CORE ;
    FOREIGN NOR3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.430 1.085 6.460 1.785 ;
        RECT  6.130 0.430 6.430 2.270 ;
        RECT  5.970 0.430 6.130 0.795 ;
        RECT  4.915 1.905 6.130 2.270 ;
        RECT  5.120 0.335 5.970 0.795 ;
        RECT  4.495 0.335 5.120 0.590 ;
        RECT  4.405 1.905 4.915 2.505 ;
        RECT  3.870 0.430 4.495 0.590 ;
        RECT  1.915 2.205 4.405 2.440 ;
        RECT  3.375 0.320 3.870 0.590 ;
        RECT  0.975 0.320 3.375 0.565 ;
        RECT  1.500 2.085 1.915 2.440 ;
        RECT  0.565 0.320 0.975 0.905 ;
        END
        AntennaDiffArea 2.381 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.720 0.975 5.950 1.440 ;
        RECT  4.940 0.975 5.720 1.135 ;
        RECT  4.780 0.770 4.940 1.135 ;
        RECT  3.295 0.770 4.780 0.930 ;
        RECT  3.195 0.770 3.295 1.345 ;
        RECT  3.035 0.745 3.195 1.345 ;
        RECT  1.320 0.745 3.035 0.905 ;
        RECT  1.160 0.745 1.320 1.245 ;
        RECT  0.720 1.085 1.160 1.245 ;
        RECT  0.560 1.085 0.720 1.580 ;
        RECT  0.390 1.225 0.560 1.580 ;
        END
        AntennaGateArea 0.7982 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.255 1.315 5.515 1.685 ;
        RECT  4.075 1.525 5.255 1.685 ;
        RECT  3.975 1.450 4.075 1.685 ;
        RECT  3.815 1.450 3.975 2.025 ;
        RECT  2.470 1.865 3.815 2.025 ;
        RECT  2.310 1.425 2.470 2.025 ;
        RECT  2.210 1.425 2.310 1.880 ;
        RECT  1.165 1.720 2.210 1.880 ;
        RECT  0.905 1.425 1.165 1.990 ;
        END
        AntennaGateArea 0.7943 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.340 1.110 4.600 1.345 ;
        RECT  3.635 1.110 4.340 1.270 ;
        RECT  3.475 1.110 3.635 1.685 ;
        RECT  2.855 1.525 3.475 1.685 ;
        RECT  2.695 1.085 2.855 1.685 ;
        RECT  2.015 1.085 2.695 1.245 ;
        RECT  1.500 1.085 2.015 1.540 ;
        END
        AntennaGateArea 0.7943 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.410 -0.130 6.560 0.130 ;
        RECT  6.150 -0.130 6.410 0.250 ;
        RECT  4.315 -0.130 6.150 0.130 ;
        RECT  4.055 -0.130 4.315 0.250 ;
        RECT  0.385 -0.130 4.055 0.130 ;
        RECT  0.125 -0.130 0.385 0.915 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.210 2.740 6.560 3.000 ;
        RECT  5.950 2.485 6.210 3.000 ;
        RECT  3.185 2.740 5.950 3.000 ;
        RECT  2.925 2.620 3.185 3.000 ;
        RECT  0.470 2.740 2.925 3.000 ;
        RECT  0.210 1.825 0.470 3.000 ;
        RECT  0.000 2.740 0.210 3.000 ;
        END
    END VDD
END NOR3X8MTH

MACRO NOR3XLMTH
    CLASS CORE ;
    FOREIGN NOR3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.710 1.950 2.035 ;
        RECT  0.615 0.710 1.740 0.920 ;
        RECT  1.505 1.795 1.740 2.035 ;
        END
        AntennaDiffArea 0.375 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.585 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 1.155 1.130 1.825 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.110 1.560 1.615 ;
        END
        AntennaGateArea 0.0702 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 -0.130 2.050 0.130 ;
        RECT  0.285 -0.130 1.225 0.390 ;
        RECT  0.000 -0.130 0.285 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.725 2.740 2.050 3.000 ;
        RECT  1.125 2.565 1.725 3.000 ;
        RECT  0.425 2.740 1.125 3.000 ;
        RECT  0.165 1.770 0.425 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
END NOR3XLMTH

MACRO NOR4BBX1MTH
    CLASS CORE ;
    FOREIGN NOR4BBX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 1.685 2.360 1.990 ;
        RECT  1.810 0.785 1.970 1.990 ;
        RECT  0.675 0.785 1.810 0.945 ;
        END
        AntennaDiffArea 0.574 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.655 1.610 ;
        END
        AntennaGateArea 0.1599 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 1.125 1.205 1.820 ;
        END
        AntennaGateArea 0.1599 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.575 1.205 3.605 1.580 ;
        RECT  3.380 0.795 3.575 1.580 ;
        END
        AntennaGateArea 0.0715 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.010 0.795 3.195 1.580 ;
        RECT  2.965 1.225 3.010 1.580 ;
        END
        AntennaGateArea 0.0715 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.390 -0.130 4.100 0.130 ;
        RECT  2.450 -0.130 3.390 0.385 ;
        RECT  1.795 -0.130 2.450 0.130 ;
        RECT  0.855 -0.130 1.795 0.385 ;
        RECT  0.385 -0.130 0.855 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.720 2.740 4.100 3.000 ;
        RECT  2.780 2.515 3.720 3.000 ;
        RECT  0.495 2.740 2.780 3.000 ;
        RECT  0.235 1.825 0.495 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.925 0.765 3.950 1.950 ;
        RECT  3.790 0.765 3.925 2.330 ;
        RECT  3.755 0.765 3.790 1.025 ;
        RECT  3.765 1.685 3.790 2.330 ;
        RECT  1.615 2.170 3.765 2.330 ;
        RECT  2.700 0.765 2.830 1.025 ;
        RECT  2.700 1.685 2.785 1.945 ;
        RECT  2.540 0.765 2.700 1.945 ;
        RECT  2.150 1.220 2.540 1.480 ;
        RECT  1.455 1.225 1.615 2.330 ;
    END
END NOR4BBX1MTH

MACRO NOR4BBX2MTH
    CLASS CORE ;
    FOREIGN NOR4BBX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.590 1.290 5.640 2.260 ;
        RECT  5.430 0.610 5.590 2.260 ;
        RECT  5.065 0.610 5.430 0.770 ;
        RECT  5.210 1.735 5.430 2.260 ;
        RECT  1.990 2.100 5.210 2.260 ;
        RECT  4.805 0.500 5.065 0.770 ;
        RECT  4.105 0.610 4.805 0.770 ;
        RECT  3.845 0.450 4.105 0.770 ;
        RECT  1.730 2.100 1.990 2.405 ;
        END
        AntennaDiffArea 1.144 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.115 0.510 3.630 0.770 ;
        END
        AntennaGateArea 0.3185 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.700 1.330 4.340 1.540 ;
        END
        AntennaGateArea 0.3185 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.160 1.350 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.450 1.075 0.730 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 0.340 ;
        RECT  3.555 -0.130 5.355 0.130 ;
        RECT  2.955 -0.130 3.555 0.275 ;
        RECT  1.035 -0.130 2.955 0.130 ;
        RECT  0.775 -0.130 1.035 0.290 ;
        RECT  0.000 -0.130 0.775 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.650 2.740 5.740 3.000 ;
        RECT  3.390 2.445 3.650 3.000 ;
        RECT  0.940 2.740 3.390 3.000 ;
        RECT  0.680 1.835 0.940 3.000 ;
        RECT  0.000 2.740 0.680 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.090 0.950 5.250 1.465 ;
        RECT  2.935 0.950 5.090 1.110 ;
        RECT  4.700 1.295 4.820 1.455 ;
        RECT  4.540 1.295 4.700 1.920 ;
        RECT  2.520 1.760 4.540 1.920 ;
        RECT  2.775 0.475 2.935 1.110 ;
        RECT  2.160 0.475 2.775 0.635 ;
        RECT  2.360 0.835 2.520 1.920 ;
        RECT  1.690 1.760 2.360 1.920 ;
        RECT  2.000 0.475 2.160 1.525 ;
        RECT  0.455 0.475 2.000 0.635 ;
        RECT  1.900 1.365 2.000 1.525 ;
        RECT  1.530 0.815 1.690 1.920 ;
        RECT  1.350 0.815 1.530 0.975 ;
        RECT  1.480 1.760 1.530 1.920 ;
        RECT  1.220 1.760 1.480 2.060 ;
        RECT  0.265 0.475 0.455 0.875 ;
        RECT  0.265 1.845 0.390 2.105 ;
        RECT  0.105 0.475 0.265 2.105 ;
    END
END NOR4BBX2MTH

MACRO NOR4BBX4MTH
    CLASS CORE ;
    FOREIGN NOR4BBX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.565 0.550 9.745 2.395 ;
        RECT  9.270 0.550 9.565 0.730 ;
        RECT  9.345 1.700 9.565 2.395 ;
        RECT  5.515 2.105 9.345 2.285 ;
        RECT  9.090 0.385 9.270 0.730 ;
        RECT  5.905 0.385 9.090 0.565 ;
        RECT  5.255 2.105 5.515 2.375 ;
        RECT  2.655 2.105 5.255 2.285 ;
        RECT  2.395 2.105 2.655 2.420 ;
        END
        AntennaDiffArea 2.024 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 1.425 7.545 1.585 ;
        RECT  3.750 1.330 4.110 1.585 ;
        END
        AntennaGateArea 0.6162 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.215 1.085 8.475 1.345 ;
        RECT  4.455 1.085 8.215 1.245 ;
        RECT  4.295 0.885 4.455 1.245 ;
        RECT  3.340 0.885 4.295 1.130 ;
        END
        AntennaGateArea 0.6162 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 1.240 1.915 1.580 ;
        END
        AntennaGateArea 0.2886 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.290 1.240 0.720 1.580 ;
        END
        AntennaGateArea 0.2886 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.715 -0.130 9.840 0.130 ;
        RECT  9.455 -0.130 9.715 0.370 ;
        RECT  5.615 -0.130 9.455 0.130 ;
        RECT  5.015 -0.130 5.615 0.520 ;
        RECT  2.545 -0.130 5.015 0.130 ;
        RECT  2.285 -0.130 2.545 0.250 ;
        RECT  1.465 -0.130 2.285 0.130 ;
        RECT  1.205 -0.130 1.465 0.250 ;
        RECT  0.385 -0.130 1.205 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.765 2.740 9.840 3.000 ;
        RECT  7.505 2.520 7.765 3.000 ;
        RECT  2.145 2.740 7.505 3.000 ;
        RECT  1.205 2.545 2.145 3.000 ;
        RECT  0.770 2.740 1.205 3.000 ;
        RECT  0.170 2.545 0.770 3.000 ;
        RECT  0.000 2.740 0.170 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.225 0.910 9.385 1.475 ;
        RECT  8.910 0.910 9.225 1.070 ;
        RECT  8.750 0.745 8.910 1.070 ;
        RECT  8.745 1.255 8.905 1.925 ;
        RECT  4.810 0.745 8.750 0.905 ;
        RECT  3.095 1.765 8.745 1.925 ;
        RECT  4.650 0.475 4.810 0.905 ;
        RECT  2.755 0.475 4.650 0.635 ;
        RECT  2.935 0.835 3.095 1.925 ;
        RECT  2.260 1.765 2.935 1.925 ;
        RECT  2.595 0.475 2.755 1.575 ;
        RECT  1.085 0.475 2.595 0.635 ;
        RECT  2.495 1.315 2.595 1.575 ;
        RECT  2.100 0.815 2.260 1.925 ;
        RECT  1.740 0.815 2.100 0.975 ;
        RECT  1.745 1.765 2.100 1.925 ;
        RECT  1.485 1.765 1.745 2.025 ;
        RECT  0.925 0.475 1.085 2.035 ;
        RECT  0.665 0.475 0.925 0.910 ;
        RECT  0.545 1.775 0.925 2.035 ;
    END
END NOR4BBX4MTH

MACRO NOR4BBXLMTH
    CLASS CORE ;
    FOREIGN NOR4BBXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.685 2.360 1.990 ;
        RECT  1.815 0.815 1.975 1.990 ;
        RECT  0.670 0.815 1.815 0.975 ;
        END
        AntennaDiffArea 0.392 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.175 0.655 1.580 ;
        END
        AntennaGateArea 0.0845 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.910 1.155 1.205 1.945 ;
        END
        AntennaGateArea 0.0845 ;
    END C
    PIN BN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.575 1.205 3.605 1.580 ;
        RECT  3.380 0.795 3.575 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END BN
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 1.225 3.195 1.930 ;
        END
        AntennaGateArea 0.0546 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.390 -0.130 4.100 0.130 ;
        RECT  2.450 -0.130 3.390 0.385 ;
        RECT  2.090 -0.130 2.450 0.130 ;
        RECT  1.490 -0.130 2.090 0.385 ;
        RECT  1.065 -0.130 1.490 0.130 ;
        RECT  0.125 -0.130 1.065 0.385 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 2.740 4.100 3.000 ;
        RECT  2.465 2.510 3.405 3.000 ;
        RECT  1.950 2.740 2.465 3.000 ;
        RECT  1.010 2.510 1.950 3.000 ;
        RECT  0.495 2.740 1.010 3.000 ;
        RECT  0.235 1.775 0.495 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.815 0.765 3.975 2.330 ;
        RECT  3.755 0.765 3.815 1.025 ;
        RECT  3.715 1.760 3.815 2.330 ;
        RECT  1.615 2.170 3.715 2.330 ;
        RECT  2.785 0.765 2.885 1.025 ;
        RECT  2.625 0.765 2.785 1.970 ;
        RECT  2.155 1.220 2.625 1.480 ;
        RECT  1.455 1.225 1.615 2.330 ;
    END
END NOR4BBXLMTH

MACRO NOR4BX1MTH
    CLASS CORE ;
    FOREIGN NOR4BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.940 2.770 2.440 ;
        RECT  2.290 0.940 2.610 1.100 ;
        RECT  2.550 1.700 2.610 2.440 ;
        RECT  2.275 1.835 2.550 2.440 ;
        RECT  2.130 0.765 2.290 1.100 ;
        RECT  1.365 0.940 2.130 1.100 ;
        RECT  1.105 0.705 1.365 1.100 ;
        END
        AntennaDiffArea 0.584 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.280 1.150 1.835 ;
        END
        AntennaGateArea 0.1599 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.280 1.755 1.795 ;
        END
        AntennaGateArea 0.1599 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 0.385 2.140 0.575 ;
        RECT  1.590 0.385 1.950 0.760 ;
        END
        AntennaGateArea 0.1599 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.045 0.355 1.625 ;
        END
        AntennaGateArea 0.0715 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 2.870 0.130 ;
        RECT  2.485 -0.130 2.745 0.415 ;
        RECT  1.375 -0.130 2.485 0.130 ;
        RECT  0.435 -0.130 1.375 0.355 ;
        RECT  0.000 -0.130 0.435 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 2.740 2.870 3.000 ;
        RECT  0.225 2.365 0.825 3.000 ;
        RECT  0.000 2.740 0.225 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.095 1.280 2.405 1.540 ;
        RECT  1.935 1.280 2.095 2.175 ;
        RECT  0.695 2.015 1.935 2.175 ;
        RECT  0.535 0.705 0.695 2.175 ;
        RECT  0.125 0.705 0.535 0.865 ;
        RECT  0.125 1.805 0.535 2.175 ;
    END
END NOR4BX1MTH

MACRO NOR4BX2MTH
    CLASS CORE ;
    FOREIGN NOR4BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.770 1.290 4.820 2.290 ;
        RECT  4.610 0.610 4.770 2.290 ;
        RECT  4.245 0.610 4.610 0.770 ;
        RECT  4.390 1.690 4.610 2.290 ;
        RECT  1.305 2.130 4.390 2.290 ;
        RECT  3.985 0.500 4.245 0.770 ;
        RECT  3.285 0.610 3.985 0.770 ;
        RECT  3.025 0.450 3.285 0.770 ;
        RECT  1.145 2.130 1.305 2.460 ;
        RECT  0.930 2.200 1.145 2.460 ;
        END
        AntennaDiffArea 1.087 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.295 0.510 2.810 0.770 ;
        END
        AntennaGateArea 0.3185 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.330 3.520 1.540 ;
        END
        AntennaGateArea 0.3185 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.880 1.295 4.000 1.455 ;
        RECT  3.720 1.295 3.880 1.900 ;
        RECT  1.990 1.740 3.720 1.900 ;
        RECT  1.720 1.740 1.990 1.950 ;
        RECT  1.560 0.835 1.720 1.950 ;
        END
        AntennaGateArea 0.3185 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.165 0.620 1.505 ;
        RECT  0.100 1.165 0.310 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.795 -0.130 4.920 0.130 ;
        RECT  4.535 -0.130 4.795 0.340 ;
        RECT  2.735 -0.130 4.535 0.130 ;
        RECT  2.135 -0.130 2.735 0.275 ;
        RECT  0.455 -0.130 2.135 0.130 ;
        RECT  0.195 -0.130 0.455 0.985 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.840 2.740 4.920 3.000 ;
        RECT  2.580 2.475 2.840 3.000 ;
        RECT  0.390 2.740 2.580 3.000 ;
        RECT  0.130 2.535 0.390 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.270 0.950 4.430 1.465 ;
        RECT  2.115 0.950 4.270 1.110 ;
        RECT  1.955 0.495 2.115 1.110 ;
        RECT  1.100 0.495 1.955 0.655 ;
        RECT  1.100 1.315 1.360 1.845 ;
        RECT  0.940 0.495 1.100 1.845 ;
        RECT  0.735 0.495 0.940 0.925 ;
        RECT  0.790 1.685 0.940 1.845 ;
        RECT  0.530 1.685 0.790 1.945 ;
    END
END NOR4BX2MTH

MACRO NOR4BX4MTH
    CLASS CORE ;
    FOREIGN NOR4BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.745 0.550 8.925 2.395 ;
        RECT  8.450 0.550 8.745 0.730 ;
        RECT  8.525 1.700 8.745 2.395 ;
        RECT  4.695 2.110 8.525 2.290 ;
        RECT  8.270 0.385 8.450 0.730 ;
        RECT  5.085 0.385 8.270 0.565 ;
        RECT  4.435 2.110 4.695 2.370 ;
        RECT  1.695 2.110 4.435 2.290 ;
        RECT  1.435 1.795 1.695 2.395 ;
        END
        AntennaDiffArea 2.02 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.325 1.425 6.725 1.585 ;
        RECT  2.725 1.330 3.325 1.585 ;
        END
        AntennaGateArea 0.6149 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.395 1.085 7.655 1.345 ;
        RECT  3.675 1.085 7.395 1.245 ;
        RECT  3.515 0.885 3.675 1.245 ;
        RECT  2.470 0.885 3.515 1.130 ;
        END
        AntennaGateArea 0.6149 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.925 1.255 8.085 1.925 ;
        RECT  2.360 1.765 7.925 1.925 ;
        RECT  2.270 1.290 2.360 1.925 ;
        RECT  1.970 0.835 2.270 1.925 ;
        END
        AntennaGateArea 0.6292 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.305 1.240 0.720 1.580 ;
        END
        AntennaGateArea 0.2886 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.895 -0.130 9.020 0.130 ;
        RECT  8.635 -0.130 8.895 0.370 ;
        RECT  4.795 -0.130 8.635 0.130 ;
        RECT  4.195 -0.130 4.795 0.520 ;
        RECT  1.415 -0.130 4.195 0.130 ;
        RECT  1.255 -0.130 1.415 1.025 ;
        RECT  0.385 -0.130 1.255 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.945 2.740 9.020 3.000 ;
        RECT  6.685 2.480 6.945 3.000 ;
        RECT  3.195 2.740 6.685 3.000 ;
        RECT  2.935 2.480 3.195 3.000 ;
        RECT  1.115 2.740 2.935 3.000 ;
        RECT  0.175 2.545 1.115 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.405 0.910 8.565 1.395 ;
        RECT  8.090 0.910 8.405 1.070 ;
        RECT  7.930 0.745 8.090 1.070 ;
        RECT  4.015 0.745 7.930 0.905 ;
        RECT  3.855 0.495 4.015 0.905 ;
        RECT  1.790 0.495 3.855 0.655 ;
        RECT  1.630 0.495 1.790 1.575 ;
        RECT  1.075 1.315 1.630 1.575 ;
        RECT  0.915 0.650 1.075 2.035 ;
        RECT  0.665 0.650 0.915 0.910 ;
        RECT  0.525 1.775 0.915 2.035 ;
    END
END NOR4BX4MTH

MACRO NOR4BXLMTH
    CLASS CORE ;
    FOREIGN NOR4BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.815 2.770 1.990 ;
        RECT  1.065 0.815 2.610 0.975 ;
        RECT  2.560 1.700 2.610 1.990 ;
        RECT  2.365 1.700 2.560 1.930 ;
        END
        AntennaDiffArea 0.392 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.155 1.150 1.755 ;
        END
        AntennaGateArea 0.0845 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.155 1.630 1.755 ;
        END
        AntennaGateArea 0.0845 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 2.110 2.360 2.435 ;
        RECT  1.715 2.275 2.150 2.435 ;
        END
        AntennaGateArea 0.0845 ;
    END B
    PIN AN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.940 0.355 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END AN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.740 -0.130 2.870 0.130 ;
        RECT  1.800 -0.130 2.740 0.380 ;
        RECT  1.260 -0.130 1.800 0.130 ;
        RECT  0.660 -0.130 1.260 0.380 ;
        RECT  0.000 -0.130 0.660 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.690 2.740 2.870 3.000 ;
        RECT  2.090 2.620 2.690 3.000 ;
        RECT  0.875 2.740 2.090 3.000 ;
        RECT  0.275 2.280 0.875 3.000 ;
        RECT  0.000 2.740 0.275 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.970 1.260 2.405 1.520 ;
        RECT  1.810 1.260 1.970 2.095 ;
        RECT  0.695 1.935 1.810 2.095 ;
        RECT  0.535 0.580 0.695 2.095 ;
        RECT  0.395 0.580 0.535 0.740 ;
        RECT  0.125 1.765 0.535 2.095 ;
        RECT  0.135 0.385 0.395 0.740 ;
    END
END NOR4BXLMTH

MACRO NOR4X12MTH
    CLASS CORE ;
    FOREIGN NOR4X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 24.190 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.480 0.310 24.020 2.440 ;
        RECT  19.395 0.310 23.480 0.530 ;
        RECT  23.265 1.495 23.480 2.440 ;
        RECT  1.665 2.145 23.265 2.440 ;
        RECT  19.110 0.310 19.395 0.590 ;
        RECT  15.860 0.430 19.110 0.590 ;
        RECT  15.530 0.310 15.860 0.590 ;
        RECT  8.290 0.310 15.530 0.565 ;
        RECT  7.915 0.310 8.290 0.590 ;
        RECT  6.950 0.430 7.915 0.590 ;
        RECT  6.590 0.310 6.950 0.590 ;
        RECT  5.495 0.310 6.590 0.565 ;
        END
        AntennaDiffArea 5.245 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.140 0.710 23.300 1.300 ;
        RECT  20.440 0.710 23.140 0.870 ;
        RECT  19.840 0.710 20.440 0.930 ;
        RECT  15.385 0.770 19.840 0.930 ;
        RECT  15.225 0.745 15.385 0.930 ;
        RECT  8.650 0.745 15.225 0.905 ;
        RECT  8.490 0.745 8.650 0.930 ;
        RECT  6.405 0.770 8.490 0.930 ;
        RECT  6.245 0.745 6.405 0.930 ;
        RECT  5.305 0.745 6.245 0.905 ;
        RECT  5.145 0.430 5.305 0.905 ;
        RECT  0.565 0.430 5.145 0.590 ;
        RECT  0.405 0.430 0.565 1.580 ;
        RECT  0.100 1.290 0.405 1.580 ;
        END
        AntennaGateArea 1.8369 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  22.410 1.050 22.870 1.210 ;
        RECT  22.250 1.050 22.410 1.955 ;
        RECT  4.115 1.795 22.250 1.955 ;
        RECT  3.855 1.450 4.115 1.955 ;
        RECT  1.130 1.795 3.855 1.955 ;
        RECT  1.105 1.290 1.130 1.955 ;
        RECT  0.745 0.835 1.105 1.955 ;
        END
        AntennaGateArea 1.8369 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.150 1.055 21.410 1.270 ;
        RECT  15.010 1.110 21.150 1.270 ;
        RECT  14.750 1.085 15.010 1.270 ;
        RECT  13.630 1.085 14.750 1.245 ;
        RECT  13.370 1.085 13.630 1.275 ;
        RECT  10.425 1.085 13.370 1.245 ;
        RECT  10.165 1.085 10.425 1.275 ;
        RECT  9.125 1.085 10.165 1.245 ;
        RECT  8.865 1.085 9.125 1.270 ;
        RECT  6.005 1.110 8.865 1.270 ;
        RECT  5.745 1.085 6.005 1.270 ;
        RECT  4.795 1.085 5.745 1.245 ;
        RECT  4.635 0.770 4.795 1.245 ;
        RECT  3.335 0.770 4.635 0.930 ;
        RECT  3.175 0.770 3.335 1.045 ;
        RECT  2.340 0.885 3.175 1.045 ;
        RECT  1.290 0.885 2.340 1.130 ;
        END
        AntennaGateArea 1.7745 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  21.680 1.315 21.840 1.615 ;
        RECT  14.340 1.455 21.680 1.615 ;
        RECT  14.080 1.425 14.340 1.615 ;
        RECT  9.795 1.455 14.080 1.615 ;
        RECT  9.535 1.425 9.795 1.615 ;
        RECT  5.255 1.455 9.535 1.615 ;
        RECT  5.045 1.425 5.255 1.615 ;
        RECT  4.455 1.425 5.045 1.585 ;
        RECT  4.295 1.110 4.455 1.585 ;
        RECT  3.675 1.110 4.295 1.270 ;
        RECT  3.515 1.110 3.675 1.575 ;
        RECT  2.095 1.415 3.515 1.575 ;
        RECT  1.495 1.330 2.095 1.575 ;
        END
        AntennaGateArea 1.7953 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.930 -0.130 24.190 0.130 ;
        RECT  18.670 -0.130 18.930 0.250 ;
        RECT  16.740 -0.130 18.670 0.130 ;
        RECT  16.140 -0.130 16.740 0.250 ;
        RECT  7.735 -0.130 16.140 0.130 ;
        RECT  7.135 -0.130 7.735 0.250 ;
        RECT  5.205 -0.130 7.135 0.130 ;
        RECT  4.945 -0.130 5.205 0.250 ;
        RECT  0.000 -0.130 4.945 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  23.740 2.740 24.190 3.000 ;
        RECT  23.140 2.620 23.740 3.000 ;
        RECT  20.400 2.740 23.140 3.000 ;
        RECT  20.140 2.620 20.400 3.000 ;
        RECT  16.550 2.740 20.140 3.000 ;
        RECT  16.290 2.620 16.550 3.000 ;
        RECT  7.585 2.740 16.290 3.000 ;
        RECT  7.325 2.620 7.585 3.000 ;
        RECT  3.425 2.740 7.325 3.000 ;
        RECT  3.165 2.620 3.425 3.000 ;
        RECT  0.455 2.740 3.165 3.000 ;
        RECT  0.195 1.835 0.455 3.000 ;
        RECT  0.000 2.740 0.195 3.000 ;
        END
    END VDD
END NOR4X12MTH

MACRO NOR4X1MTH
    CLASS CORE ;
    FOREIGN NOR4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.805 2.370 2.460 ;
        RECT  1.905 0.805 2.210 0.965 ;
        RECT  2.150 1.700 2.210 2.460 ;
        RECT  1.990 1.860 2.150 2.460 ;
        RECT  1.645 0.705 1.905 0.965 ;
        RECT  0.905 0.805 1.645 0.965 ;
        RECT  0.645 0.705 0.905 0.965 ;
        END
        AntennaDiffArea 0.574 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.155 0.600 1.520 ;
        RECT  0.100 1.155 0.310 1.665 ;
        END
        AntennaGateArea 0.1599 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.820 1.280 1.080 1.990 ;
        RECT  0.510 1.700 0.820 1.990 ;
        END
        AntennaGateArea 0.1599 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 1.225 1.550 1.845 ;
        END
        AntennaGateArea 0.1599 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.145 2.030 1.485 ;
        RECT  1.730 1.145 1.950 1.680 ;
        END
        AntennaGateArea 0.1599 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  1.395 -0.130 2.335 0.355 ;
        RECT  1.070 -0.130 1.395 0.130 ;
        RECT  0.390 -0.130 1.070 0.355 ;
        RECT  0.130 -0.130 0.390 0.965 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.390 2.740 2.460 3.000 ;
        RECT  0.130 2.170 0.390 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
END NOR4X1MTH

MACRO NOR4X2MTH
    CLASS CORE ;
    FOREIGN NOR4X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.950 1.290 4.000 1.800 ;
        RECT  3.790 0.610 3.950 1.800 ;
        RECT  3.425 0.610 3.790 0.770 ;
        RECT  3.400 1.640 3.790 1.800 ;
        RECT  3.165 0.500 3.425 0.770 ;
        RECT  3.240 1.640 3.400 2.290 ;
        RECT  2.050 2.130 3.240 2.290 ;
        RECT  2.465 0.610 3.165 0.770 ;
        RECT  2.205 0.450 2.465 0.770 ;
        RECT  1.790 2.130 2.050 2.395 ;
        END
        AntennaDiffArea 0.894 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 0.950 3.610 1.455 ;
        RECT  1.305 0.950 3.450 1.110 ;
        RECT  1.145 0.495 1.305 1.110 ;
        RECT  0.535 0.495 1.145 0.655 ;
        RECT  0.375 0.495 0.535 1.580 ;
        RECT  0.100 1.260 0.375 1.580 ;
        END
        AntennaGateArea 0.3185 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.060 1.295 3.180 1.455 ;
        RECT  2.900 1.295 3.060 1.900 ;
        RECT  1.170 1.740 2.900 1.900 ;
        RECT  0.945 1.740 1.170 1.950 ;
        RECT  0.785 0.835 0.945 1.950 ;
        END
        AntennaGateArea 0.3185 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.125 1.330 2.700 1.540 ;
        END
        AntennaGateArea 0.3185 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.485 0.510 1.990 0.770 ;
        END
        AntennaGateArea 0.3185 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.100 0.130 ;
        RECT  3.715 -0.130 3.975 0.340 ;
        RECT  1.925 -0.130 3.715 0.130 ;
        RECT  1.325 -0.130 1.925 0.275 ;
        RECT  0.000 -0.130 1.325 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.870 2.740 4.100 3.000 ;
        RECT  3.610 1.980 3.870 3.000 ;
        RECT  0.410 2.740 3.610 3.000 ;
        RECT  0.150 1.875 0.410 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
END NOR4X2MTH

MACRO NOR4X4MTH
    CLASS CORE ;
    FOREIGN NOR4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.515 0.595 7.695 1.760 ;
        RECT  7.220 0.595 7.515 0.775 ;
        RECT  7.215 1.580 7.515 1.760 ;
        RECT  7.040 0.375 7.220 0.775 ;
        RECT  7.035 1.580 7.215 2.285 ;
        RECT  3.855 0.375 7.040 0.565 ;
        RECT  5.735 2.105 7.035 2.285 ;
        RECT  5.430 2.105 5.735 2.400 ;
        RECT  1.925 2.105 5.430 2.285 ;
        RECT  1.665 2.105 1.925 2.390 ;
        END
        AntennaDiffArea 1.849 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.175 0.960 7.335 1.395 ;
        RECT  6.815 0.960 7.175 1.120 ;
        RECT  6.655 0.745 6.815 1.120 ;
        RECT  3.115 0.745 6.655 0.905 ;
        RECT  2.955 0.495 3.115 0.905 ;
        RECT  0.560 0.495 2.955 0.655 ;
        RECT  0.400 0.495 0.560 1.580 ;
        RECT  0.100 1.290 0.400 1.580 ;
        END
        AntennaGateArea 0.637 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.695 1.315 6.855 1.925 ;
        RECT  1.130 1.765 6.695 1.925 ;
        RECT  1.060 1.290 1.130 1.925 ;
        RECT  0.740 0.835 1.060 1.925 ;
        END
        AntennaGateArea 0.6292 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.165 1.085 6.425 1.345 ;
        RECT  2.450 1.085 6.165 1.245 ;
        RECT  2.290 0.885 2.450 1.245 ;
        RECT  1.290 0.885 2.290 1.130 ;
        END
        AntennaGateArea 0.6149 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.095 1.425 5.480 1.585 ;
        RECT  1.495 1.330 2.095 1.585 ;
        END
        AntennaGateArea 0.6149 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 -0.130 7.790 0.130 ;
        RECT  7.405 -0.130 7.665 0.375 ;
        RECT  3.595 -0.130 7.405 0.130 ;
        RECT  3.335 -0.130 3.595 0.565 ;
        RECT  0.000 -0.130 3.335 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.570 2.740 7.790 3.000 ;
        RECT  7.410 1.985 7.570 3.000 ;
        RECT  3.425 2.740 7.410 3.000 ;
        RECT  3.165 2.505 3.425 3.000 ;
        RECT  0.460 2.740 3.165 3.000 ;
        RECT  0.200 1.835 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
END NOR4X4MTH

MACRO NOR4X6MTH
    CLASS CORE ;
    FOREIGN NOR4X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.555 0.615 11.800 2.410 ;
        RECT  11.325 0.615 11.555 0.905 ;
        RECT  1.665 2.130 11.555 2.410 ;
        RECT  10.955 0.310 11.325 0.905 ;
        RECT  8.290 0.310 10.955 0.565 ;
        RECT  7.915 0.310 8.290 0.590 ;
        RECT  6.955 0.430 7.915 0.590 ;
        RECT  6.680 0.310 6.955 0.590 ;
        RECT  5.495 0.310 6.680 0.565 ;
        END
        AntennaDiffArea 2.771 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.215 1.085 11.375 1.460 ;
        RECT  10.775 1.085 11.215 1.245 ;
        RECT  10.615 0.745 10.775 1.245 ;
        RECT  8.650 0.745 10.615 0.905 ;
        RECT  8.490 0.745 8.650 0.930 ;
        RECT  6.405 0.770 8.490 0.930 ;
        RECT  6.245 0.745 6.405 0.930 ;
        RECT  5.305 0.745 6.245 0.905 ;
        RECT  5.145 0.430 5.305 0.905 ;
        RECT  0.560 0.430 5.145 0.590 ;
        RECT  0.400 0.430 0.560 1.580 ;
        RECT  0.100 1.290 0.400 1.580 ;
        END
        AntennaGateArea 0.936 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 1.425 10.945 1.585 ;
        RECT  10.685 1.425 10.845 1.950 ;
        RECT  4.115 1.790 10.685 1.950 ;
        RECT  3.855 1.450 4.115 1.950 ;
        RECT  1.130 1.790 3.855 1.950 ;
        RECT  1.105 1.290 1.130 1.950 ;
        RECT  0.740 0.835 1.105 1.950 ;
        END
        AntennaGateArea 0.9217 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.365 1.355 10.465 1.515 ;
        RECT  10.205 1.085 10.365 1.515 ;
        RECT  9.125 1.085 10.205 1.245 ;
        RECT  8.865 1.085 9.125 1.270 ;
        RECT  6.005 1.110 8.865 1.270 ;
        RECT  5.745 1.085 6.005 1.270 ;
        RECT  4.795 1.085 5.745 1.245 ;
        RECT  4.635 0.770 4.795 1.245 ;
        RECT  3.335 0.770 4.635 0.930 ;
        RECT  3.175 0.770 3.335 1.045 ;
        RECT  2.340 0.885 3.175 1.045 ;
        RECT  1.290 0.885 2.340 1.130 ;
        END
        AntennaGateArea 0.9009 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.385 1.425 9.985 1.610 ;
        RECT  5.255 1.450 9.385 1.610 ;
        RECT  5.045 1.425 5.255 1.610 ;
        RECT  4.455 1.425 5.045 1.585 ;
        RECT  4.295 1.110 4.455 1.585 ;
        RECT  3.675 1.110 4.295 1.270 ;
        RECT  3.515 1.110 3.675 1.575 ;
        RECT  2.095 1.415 3.515 1.575 ;
        RECT  1.495 1.330 2.095 1.575 ;
        END
        AntennaGateArea 0.9113 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 -0.130 11.890 0.130 ;
        RECT  11.505 -0.130 11.765 0.300 ;
        RECT  7.735 -0.130 11.505 0.130 ;
        RECT  7.135 -0.130 7.735 0.250 ;
        RECT  5.205 -0.130 7.135 0.130 ;
        RECT  4.945 -0.130 5.205 0.250 ;
        RECT  0.000 -0.130 4.945 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.625 2.740 11.890 3.000 ;
        RECT  11.365 2.620 11.625 3.000 ;
        RECT  7.585 2.740 11.365 3.000 ;
        RECT  7.325 2.590 7.585 3.000 ;
        RECT  3.425 2.740 7.325 3.000 ;
        RECT  3.165 2.620 3.425 3.000 ;
        RECT  0.460 2.740 3.165 3.000 ;
        RECT  0.200 1.835 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
END NOR4X6MTH

MACRO NOR4X8MTH
    CLASS CORE ;
    FOREIGN NOR4X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.990 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.385 0.310 15.785 2.440 ;
        RECT  12.755 0.310 15.385 0.590 ;
        RECT  15.270 1.475 15.385 2.440 ;
        RECT  1.665 2.170 15.270 2.440 ;
        RECT  12.135 0.430 12.755 0.590 ;
        RECT  11.750 0.310 12.135 0.590 ;
        RECT  8.765 0.310 11.750 0.565 ;
        RECT  8.325 0.310 8.765 0.590 ;
        RECT  7.265 0.430 8.325 0.590 ;
        RECT  7.010 0.310 7.265 0.590 ;
        RECT  3.855 0.310 7.010 0.565 ;
        END
        AntennaDiffArea 3.604 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.500 0.770 12.940 0.930 ;
        RECT  11.340 0.745 11.500 0.930 ;
        RECT  9.150 0.745 11.340 0.905 ;
        RECT  8.990 0.745 9.150 0.930 ;
        RECT  6.815 0.770 8.990 0.930 ;
        RECT  6.655 0.745 6.815 0.930 ;
        RECT  3.115 0.745 6.655 0.905 ;
        RECT  2.955 0.495 3.115 0.905 ;
        RECT  0.565 0.495 2.955 0.655 ;
        RECT  0.405 0.495 0.565 1.580 ;
        RECT  0.100 1.290 0.405 1.580 ;
        END
        AntennaGateArea 1.274 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.015 0.905 15.205 1.165 ;
        RECT  14.855 0.905 15.015 1.950 ;
        RECT  1.130 1.790 14.855 1.950 ;
        RECT  1.105 1.290 1.130 1.950 ;
        RECT  0.745 0.835 1.105 1.950 ;
        END
        AntennaGateArea 1.2428 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.485 0.980 13.745 1.270 ;
        RECT  11.145 1.110 13.485 1.270 ;
        RECT  11.025 1.085 11.145 1.270 ;
        RECT  9.745 1.085 11.025 1.245 ;
        RECT  9.550 1.085 9.745 1.270 ;
        RECT  6.425 1.110 9.550 1.270 ;
        RECT  6.160 1.085 6.425 1.270 ;
        RECT  2.450 1.085 6.160 1.245 ;
        RECT  2.290 0.885 2.450 1.245 ;
        RECT  1.290 0.885 2.290 1.130 ;
        END
        AntennaGateArea 1.1934 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.145 1.315 14.405 1.610 ;
        RECT  10.590 1.450 14.145 1.610 ;
        RECT  9.990 1.425 10.590 1.610 ;
        RECT  5.815 1.450 9.990 1.610 ;
        RECT  5.575 1.425 5.815 1.610 ;
        RECT  2.095 1.425 5.575 1.585 ;
        RECT  1.495 1.330 2.095 1.585 ;
        END
        AntennaGateArea 1.2142 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.570 -0.130 15.990 0.130 ;
        RECT  12.310 -0.130 12.570 0.250 ;
        RECT  8.145 -0.130 12.310 0.130 ;
        RECT  7.545 -0.130 8.145 0.250 ;
        RECT  3.595 -0.130 7.545 0.130 ;
        RECT  3.335 -0.130 3.595 0.565 ;
        RECT  0.000 -0.130 3.335 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.735 2.740 15.990 3.000 ;
        RECT  15.475 2.620 15.735 3.000 ;
        RECT  12.715 2.740 15.475 3.000 ;
        RECT  12.455 2.620 12.715 3.000 ;
        RECT  7.995 2.740 12.455 3.000 ;
        RECT  7.735 2.620 7.995 3.000 ;
        RECT  3.425 2.740 7.735 3.000 ;
        RECT  3.165 2.620 3.425 3.000 ;
        RECT  0.460 2.740 3.165 3.000 ;
        RECT  0.200 1.835 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
END NOR4X8MTH

MACRO NOR4XLMTH
    CLASS CORE ;
    FOREIGN NOR4XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.805 2.360 2.135 ;
        RECT  1.885 0.805 2.200 0.965 ;
        RECT  2.150 1.700 2.200 2.135 ;
        RECT  1.990 1.905 2.150 2.135 ;
        RECT  1.625 0.705 1.885 0.965 ;
        RECT  0.845 0.805 1.625 0.965 ;
        RECT  0.585 0.705 0.845 0.965 ;
        END
        AntennaDiffArea 0.43 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.155 0.600 1.520 ;
        RECT  0.100 1.155 0.310 1.855 ;
        END
        AntennaGateArea 0.0845 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 1.280 1.085 1.990 ;
        RECT  0.510 1.700 0.825 1.990 ;
        END
        AntennaGateArea 0.0845 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.270 1.225 1.550 1.845 ;
        END
        AntennaGateArea 0.0845 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.145 2.020 1.485 ;
        RECT  1.730 1.145 1.950 1.680 ;
        END
        AntennaGateArea 0.0845 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  1.395 -0.130 2.335 0.445 ;
        RECT  1.065 -0.130 1.395 0.130 ;
        RECT  0.125 -0.130 1.065 0.445 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 2.740 2.460 3.000 ;
        RECT  1.010 2.565 1.950 3.000 ;
        RECT  0.385 2.740 1.010 3.000 ;
        RECT  0.125 2.170 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END NOR4XLMTH

MACRO OA21X1MTH
    CLASS CORE ;
    FOREIGN OA21X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 1.290 2.770 1.580 ;
        RECT  2.720 0.415 2.745 0.675 ;
        RECT  2.720 1.940 2.745 2.200 ;
        RECT  2.560 0.415 2.720 2.200 ;
        RECT  2.485 0.415 2.560 0.675 ;
        RECT  2.485 1.940 2.560 2.200 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.205 1.655 1.655 ;
        END
        AntennaGateArea 0.0598 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.595 1.610 ;
        END
        AntennaGateArea 0.0598 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.775 1.205 1.130 1.655 ;
        END
        AntennaGateArea 0.0598 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 -0.130 2.870 0.130 ;
        RECT  1.945 -0.130 2.205 0.675 ;
        RECT  1.545 -0.130 1.945 0.130 ;
        RECT  1.285 -0.130 1.545 0.340 ;
        RECT  0.965 -0.130 1.285 0.130 ;
        RECT  0.705 -0.130 0.965 0.685 ;
        RECT  0.000 -0.130 0.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.185 2.740 2.870 3.000 ;
        RECT  1.585 2.225 2.185 3.000 ;
        RECT  1.335 2.740 1.585 3.000 ;
        RECT  0.735 2.485 1.335 3.000 ;
        RECT  0.385 2.740 0.735 3.000 ;
        RECT  0.125 1.845 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.115 1.315 2.380 1.575 ;
        RECT  1.955 0.925 2.115 1.995 ;
        RECT  1.855 0.925 1.955 1.185 ;
        RECT  1.275 1.835 1.955 1.995 ;
        RECT  1.285 0.765 1.545 1.025 ;
        RECT  0.385 0.865 1.285 1.025 ;
        RECT  1.015 1.835 1.275 2.105 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END OA21X1MTH

MACRO OA21X2MTH
    CLASS CORE ;
    FOREIGN OA21X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 1.700 2.770 2.410 ;
        RECT  2.695 0.380 2.745 0.980 ;
        RECT  2.535 0.380 2.695 2.410 ;
        RECT  2.485 0.380 2.535 0.980 ;
        RECT  2.475 1.700 2.535 2.410 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.185 1.630 1.580 ;
        END
        AntennaGateArea 0.0949 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.330 1.135 0.355 1.520 ;
        RECT  0.100 1.135 0.330 1.910 ;
        END
        AntennaGateArea 0.0949 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.025 1.225 1.075 1.485 ;
        RECT  0.815 1.225 1.025 1.580 ;
        RECT  0.720 1.420 0.815 1.580 ;
        RECT  0.560 1.420 0.720 1.990 ;
        RECT  0.510 1.700 0.560 1.990 ;
        END
        AntennaGateArea 0.0949 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.205 -0.130 2.870 0.130 ;
        RECT  1.605 -0.130 2.205 0.460 ;
        RECT  0.855 -0.130 1.605 0.130 ;
        RECT  0.595 -0.130 0.855 0.975 ;
        RECT  0.000 -0.130 0.595 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 2.740 2.870 3.000 ;
        RECT  1.580 2.230 2.180 3.000 ;
        RECT  0.385 2.740 1.580 3.000 ;
        RECT  0.125 2.185 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.145 1.185 2.355 1.445 ;
        RECT  1.985 0.835 2.145 1.920 ;
        RECT  1.795 0.835 1.985 0.995 ;
        RECT  1.245 1.760 1.985 1.920 ;
        RECT  1.535 0.735 1.795 0.995 ;
        RECT  0.985 1.760 1.245 2.035 ;
    END
END OA21X2MTH

MACRO OA21X4MTH
    CLASS CORE ;
    FOREIGN OA21X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 0.380 3.055 0.980 ;
        RECT  2.795 0.380 2.975 1.870 ;
        RECT  2.360 1.690 2.795 1.870 ;
        RECT  2.150 1.690 2.360 2.410 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.160 1.630 1.595 ;
        END
        AntennaGateArea 0.1885 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.600 1.660 ;
        END
        AntennaGateArea 0.1885 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 0.880 1.130 1.485 ;
        RECT  0.855 1.225 0.920 1.485 ;
        END
        AntennaGateArea 0.1885 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.560 -0.130 3.690 0.130 ;
        RECT  3.310 -0.130 3.560 0.980 ;
        RECT  2.545 -0.130 3.310 0.130 ;
        RECT  2.285 -0.130 2.545 0.980 ;
        RECT  0.935 -0.130 2.285 0.130 ;
        RECT  0.675 -0.130 0.935 0.335 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.260 2.740 3.690 3.000 ;
        RECT  2.660 2.230 3.260 3.000 ;
        RECT  1.840 2.740 2.660 3.000 ;
        RECT  1.580 2.230 1.840 3.000 ;
        RECT  0.425 2.740 1.580 3.000 ;
        RECT  0.165 1.865 0.425 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.970 1.205 2.615 1.465 ;
        RECT  1.970 0.380 1.995 0.980 ;
        RECT  1.810 0.380 1.970 1.935 ;
        RECT  1.735 0.380 1.810 0.980 ;
        RECT  1.285 1.775 1.810 1.935 ;
        RECT  1.225 0.440 1.485 0.700 ;
        RECT  1.025 1.775 1.285 2.375 ;
        RECT  0.390 0.540 1.225 0.700 ;
        RECT  0.130 0.380 0.390 0.980 ;
    END
END OA21X4MTH

MACRO OA21X8MTH
    CLASS CORE ;
    FOREIGN OA21X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.620 0.380 5.970 2.390 ;
        RECT  5.430 0.880 5.620 1.785 ;
        RECT  5.055 1.180 5.430 1.530 ;
        RECT  4.705 0.380 5.055 2.410 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.225 3.625 1.580 ;
        END
        AntennaGateArea 0.377 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.225 1.065 1.580 ;
        END
        AntennaGateArea 0.377 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.225 2.060 1.580 ;
        END
        AntennaGateArea 0.377 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.980 ;
        RECT  2.450 -0.130 6.175 0.130 ;
        RECT  2.190 -0.130 2.450 0.635 ;
        RECT  1.425 -0.130 2.190 0.130 ;
        RECT  1.165 -0.130 1.425 0.635 ;
        RECT  0.385 -0.130 1.165 0.130 ;
        RECT  0.125 -0.130 0.385 0.985 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.385 2.740 6.560 3.000 ;
        RECT  6.185 1.790 6.385 3.000 ;
        RECT  4.425 2.740 6.185 3.000 ;
        RECT  4.165 2.570 4.425 3.000 ;
        RECT  3.485 2.740 4.165 3.000 ;
        RECT  3.225 2.105 3.485 3.000 ;
        RECT  0.905 2.740 3.225 3.000 ;
        RECT  0.645 2.105 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.965 1.230 4.525 1.490 ;
        RECT  3.735 0.355 3.995 0.615 ;
        RECT  3.965 1.760 3.995 2.315 ;
        RECT  3.805 0.845 3.965 2.315 ;
        RECT  3.485 0.845 3.805 1.005 ;
        RECT  3.735 1.760 3.805 2.315 ;
        RECT  2.975 0.405 3.735 0.565 ;
        RECT  2.975 1.760 3.735 1.920 ;
        RECT  3.225 0.745 3.485 1.005 ;
        RECT  2.715 0.375 2.975 0.975 ;
        RECT  2.715 1.760 2.975 2.360 ;
        RECT  1.935 0.815 2.715 0.975 ;
        RECT  1.935 1.760 2.715 1.920 ;
        RECT  2.185 2.125 2.445 2.360 ;
        RECT  1.425 2.200 2.185 2.360 ;
        RECT  1.675 0.375 1.935 0.975 ;
        RECT  1.675 1.760 1.935 2.020 ;
        RECT  0.905 0.815 1.675 0.975 ;
        RECT  1.165 1.760 1.425 2.360 ;
        RECT  0.385 1.760 1.165 1.920 ;
        RECT  0.645 0.375 0.905 0.975 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END OA21X8MTH

MACRO OA21XLMTH
    CLASS CORE ;
    FOREIGN OA21XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 1.290 2.770 1.580 ;
        RECT  2.720 0.525 2.745 0.785 ;
        RECT  2.720 1.835 2.745 2.095 ;
        RECT  2.560 0.525 2.720 2.095 ;
        RECT  2.485 0.525 2.560 0.785 ;
        RECT  2.485 1.835 2.560 2.095 ;
        END
        AntennaDiffArea 0.236 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.205 1.655 1.655 ;
        END
        AntennaGateArea 0.0598 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.595 1.610 ;
        END
        AntennaGateArea 0.0598 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.775 1.205 1.130 1.655 ;
        END
        AntennaGateArea 0.0598 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 -0.130 2.870 0.130 ;
        RECT  1.915 -0.130 2.175 0.665 ;
        RECT  1.535 -0.130 1.915 0.130 ;
        RECT  1.275 -0.130 1.535 0.355 ;
        RECT  0.965 -0.130 1.275 0.130 ;
        RECT  0.705 -0.130 0.965 0.685 ;
        RECT  0.000 -0.130 0.705 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 2.740 2.870 3.000 ;
        RECT  1.575 2.345 2.175 3.000 ;
        RECT  1.300 2.740 1.575 3.000 ;
        RECT  0.700 2.345 1.300 3.000 ;
        RECT  0.385 2.740 0.700 3.000 ;
        RECT  0.125 1.835 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.115 1.305 2.375 1.565 ;
        RECT  1.955 0.915 2.115 1.995 ;
        RECT  1.855 0.915 1.955 1.175 ;
        RECT  1.275 1.835 1.955 1.995 ;
        RECT  1.285 0.765 1.545 1.025 ;
        RECT  0.385 0.865 1.285 1.025 ;
        RECT  1.015 1.835 1.275 2.095 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END OA21XLMTH

MACRO OA22X1MTH
    CLASS CORE ;
    FOREIGN OA22X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 0.740 3.180 2.115 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 1.245 2.360 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 1.115 1.645 1.610 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.370 1.245 0.445 1.505 ;
        RECT  0.100 0.880 0.370 1.505 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 2.190 1.075 2.350 ;
        RECT  0.565 1.700 0.725 2.350 ;
        RECT  0.510 1.700 0.565 1.990 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 -0.130 3.280 0.130 ;
        RECT  2.805 -0.130 3.065 0.290 ;
        RECT  2.555 -0.130 2.805 0.130 ;
        RECT  1.615 -0.130 2.555 0.385 ;
        RECT  0.000 -0.130 1.615 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.590 2.740 3.280 3.000 ;
        RECT  2.330 2.150 2.590 3.000 ;
        RECT  1.685 2.740 2.330 3.000 ;
        RECT  0.745 2.585 1.685 3.000 ;
        RECT  0.385 2.740 0.745 3.000 ;
        RECT  0.125 2.180 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.555 1.285 2.715 1.970 ;
        RECT  1.120 1.810 2.555 1.970 ;
        RECT  1.985 0.765 2.245 1.045 ;
        RECT  1.305 0.765 1.985 0.925 ;
        RECT  1.145 0.355 1.305 0.925 ;
        RECT  1.045 0.355 1.145 0.515 ;
        RECT  0.960 1.310 1.120 1.970 ;
        RECT  0.815 1.310 0.960 1.470 ;
        RECT  0.655 0.765 0.815 1.470 ;
        RECT  0.555 0.765 0.655 1.025 ;
    END
END OA22X1MTH

MACRO OA22X2MTH
    CLASS CORE ;
    FOREIGN OA22X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 0.410 3.180 2.380 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.820 1.205 2.360 1.580 ;
        END
        AntennaGateArea 0.1131 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.240 1.210 1.630 1.580 ;
        END
        AntennaGateArea 0.1131 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 0.565 1.520 ;
        RECT  0.100 1.205 0.310 1.580 ;
        END
        AntennaGateArea 0.1131 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 2.315 1.210 2.475 ;
        RECT  0.560 1.700 0.720 2.475 ;
        RECT  0.510 1.700 0.560 1.990 ;
        END
        AntennaGateArea 0.1131 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 -0.130 3.280 0.130 ;
        RECT  1.620 -0.130 2.560 0.415 ;
        RECT  0.000 -0.130 1.620 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.580 2.740 3.280 3.000 ;
        RECT  1.980 2.140 2.580 3.000 ;
        RECT  0.380 2.740 1.980 3.000 ;
        RECT  0.220 2.180 0.380 3.000 ;
        RECT  0.000 2.740 0.220 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.555 1.255 2.715 1.920 ;
        RECT  1.380 1.760 2.555 1.920 ;
        RECT  1.085 0.765 2.245 1.025 ;
        RECT  1.120 1.760 1.380 2.020 ;
        RECT  1.060 1.760 1.120 1.920 ;
        RECT  0.905 1.205 1.060 1.920 ;
        RECT  0.900 0.765 0.905 1.920 ;
        RECT  0.745 0.765 0.900 1.365 ;
        RECT  0.525 0.765 0.745 1.025 ;
    END
END OA22X2MTH

MACRO OA22X4MTH
    CLASS CORE ;
    FOREIGN OA22X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 1.205 3.590 1.580 ;
        RECT  3.205 0.400 3.465 2.375 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.190 2.610 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.155 1.630 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.565 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.155 1.130 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.100 0.130 ;
        RECT  3.715 -0.130 3.975 1.000 ;
        RECT  2.955 -0.130 3.715 0.130 ;
        RECT  2.695 -0.130 2.955 0.985 ;
        RECT  0.000 -0.130 2.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 1.785 3.975 3.000 ;
        RECT  2.865 2.740 3.715 3.000 ;
        RECT  2.265 2.110 2.865 3.000 ;
        RECT  0.385 2.740 2.265 3.000 ;
        RECT  0.125 1.845 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.865 1.230 3.025 1.930 ;
        RECT  1.970 1.770 2.865 1.930 ;
        RECT  2.180 0.405 2.440 1.005 ;
        RECT  0.385 0.405 2.180 0.565 ;
        RECT  1.810 0.815 1.970 1.930 ;
        RECT  0.635 0.815 1.810 0.975 ;
        RECT  1.555 1.770 1.810 1.930 ;
        RECT  0.955 1.770 1.555 2.415 ;
        RECT  0.125 0.405 0.385 1.005 ;
    END
END OA22X4MTH

MACRO OA22X8MTH
    CLASS CORE ;
    FOREIGN OA22X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.030 0.400 6.380 2.375 ;
        RECT  5.415 1.290 6.030 1.575 ;
        RECT  5.065 0.400 5.415 2.375 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.890 1.290 3.525 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 1.290 4.125 1.580 ;
        RECT  3.705 1.290 3.865 1.920 ;
        RECT  2.695 1.760 3.705 1.920 ;
        RECT  2.535 1.245 2.695 1.920 ;
        RECT  2.345 1.245 2.535 1.505 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.250 1.540 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 1.275 2.125 1.535 ;
        RECT  1.855 1.275 2.015 1.880 ;
        RECT  0.505 1.720 1.855 1.880 ;
        RECT  0.100 1.235 0.505 1.880 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 -0.130 6.970 0.130 ;
        RECT  6.585 -0.130 6.845 0.980 ;
        RECT  5.800 -0.130 6.585 0.130 ;
        RECT  5.595 -0.130 5.800 1.000 ;
        RECT  4.775 -0.130 5.595 0.130 ;
        RECT  4.515 -0.130 4.775 0.295 ;
        RECT  0.000 -0.130 4.515 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 1.785 6.845 3.000 ;
        RECT  5.775 2.740 6.585 3.000 ;
        RECT  5.595 1.785 5.775 3.000 ;
        RECT  4.765 2.740 5.595 3.000 ;
        RECT  4.505 2.100 4.765 3.000 ;
        RECT  3.340 2.740 4.505 3.000 ;
        RECT  3.080 2.440 3.340 3.000 ;
        RECT  1.310 2.740 3.080 3.000 ;
        RECT  1.050 2.440 1.310 3.000 ;
        RECT  0.000 2.740 1.050 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.545 1.230 4.885 1.490 ;
        RECT  4.385 0.950 4.545 1.920 ;
        RECT  3.055 0.950 4.385 1.110 ;
        RECT  4.245 1.760 4.385 1.920 ;
        RECT  3.415 0.610 4.365 0.770 ;
        RECT  4.045 1.760 4.245 2.360 ;
        RECT  2.355 2.100 4.045 2.260 ;
        RECT  3.255 0.405 3.415 0.770 ;
        RECT  0.385 0.405 3.255 0.565 ;
        RECT  2.895 0.815 3.055 1.110 ;
        RECT  0.635 0.815 2.895 0.975 ;
        RECT  2.195 1.800 2.355 2.400 ;
        RECT  0.385 2.100 2.195 2.260 ;
        RECT  0.125 0.405 0.385 1.005 ;
        RECT  0.125 2.100 0.385 2.360 ;
    END
END OA22X8MTH

MACRO OA22XLMTH
    CLASS CORE ;
    FOREIGN OA22XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.895 0.335 3.180 2.115 ;
        END
        AntennaDiffArea 0.337 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 1.245 2.360 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 1.115 1.645 1.610 ;
        END
        AntennaGateArea 0.0533 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.370 1.245 0.445 1.505 ;
        RECT  0.100 0.880 0.370 1.505 ;
        END
        AntennaGateArea 0.0533 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 2.160 1.075 2.320 ;
        RECT  0.565 1.700 0.725 2.320 ;
        RECT  0.510 1.700 0.565 1.990 ;
        END
        AntennaGateArea 0.0533 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.555 -0.130 3.280 0.130 ;
        RECT  1.615 -0.130 2.555 0.385 ;
        RECT  0.000 -0.130 1.615 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.590 2.740 3.280 3.000 ;
        RECT  2.330 2.140 2.590 3.000 ;
        RECT  1.685 2.740 2.330 3.000 ;
        RECT  0.745 2.585 1.685 3.000 ;
        RECT  0.385 2.740 0.745 3.000 ;
        RECT  0.125 2.180 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.555 1.285 2.715 1.950 ;
        RECT  1.120 1.790 2.555 1.950 ;
        RECT  1.985 0.765 2.245 1.025 ;
        RECT  1.305 0.765 1.985 0.925 ;
        RECT  1.145 0.385 1.305 0.925 ;
        RECT  1.045 0.385 1.145 0.545 ;
        RECT  0.960 1.310 1.120 1.950 ;
        RECT  0.815 1.310 0.960 1.470 ;
        RECT  0.655 0.765 0.815 1.470 ;
        RECT  0.555 0.765 0.655 1.025 ;
    END
END OA22XLMTH

MACRO OAI211X1MTH
    CLASS CORE ;
    FOREIGN OAI211X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 0.770 2.370 1.990 ;
        RECT  1.990 0.770 2.210 0.930 ;
        RECT  2.150 1.700 2.210 1.990 ;
        RECT  1.275 1.830 2.150 1.990 ;
        RECT  1.115 1.830 1.275 2.330 ;
        RECT  0.335 2.170 1.115 2.330 ;
        RECT  0.175 2.070 0.335 2.330 ;
        END
        AntennaDiffArea 0.581 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 1.175 1.550 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.110 2.030 1.540 ;
        RECT  1.730 1.110 1.990 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.760 1.315 1.005 1.575 ;
        RECT  0.535 1.315 0.760 1.950 ;
        RECT  0.470 1.740 0.535 1.950 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.120 0.355 1.600 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 -0.130 2.460 0.130 ;
        RECT  1.575 -0.130 2.175 0.405 ;
        RECT  1.275 -0.130 1.575 0.130 ;
        RECT  0.675 -0.130 1.275 0.405 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  2.075 2.170 2.335 3.000 ;
        RECT  1.235 2.740 2.075 3.000 ;
        RECT  0.975 2.510 1.235 3.000 ;
        RECT  0.000 2.740 0.975 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.125 0.780 1.420 0.940 ;
    END
END OAI211X1MTH

MACRO OAI211X2MTH
    CLASS CORE ;
    FOREIGN OAI211X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.045 0.355 2.305 0.955 ;
        RECT  1.900 0.470 2.045 0.955 ;
        RECT  1.740 0.470 1.900 2.330 ;
        RECT  0.395 2.170 1.740 2.330 ;
        RECT  0.135 2.170 0.395 2.430 ;
        END
        AntennaDiffArea 0.871 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.215 1.540 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.080 1.215 2.360 1.855 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.700 1.215 1.000 1.990 ;
        RECT  0.470 1.740 0.700 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.135 0.515 1.560 ;
        RECT  0.100 1.135 0.310 1.640 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 -0.130 2.460 0.130 ;
        RECT  0.645 -0.130 0.905 0.615 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.320 2.740 2.460 3.000 ;
        RECT  2.110 2.035 2.320 3.000 ;
        RECT  0.000 2.740 2.110 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.195 0.355 1.455 0.955 ;
        RECT  0.385 0.795 1.195 0.955 ;
        RECT  0.125 0.355 0.385 0.955 ;
    END
END OAI211X2MTH

MACRO OAI211X4MTH
    CLASS CORE ;
    FOREIGN OAI211X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.365 1.290 4.410 1.580 ;
        RECT  4.105 0.745 4.365 2.310 ;
        RECT  3.005 0.745 4.105 0.905 ;
        RECT  2.165 2.130 4.105 2.310 ;
        RECT  1.905 1.955 2.165 2.455 ;
        RECT  0.445 1.955 1.905 2.135 ;
        RECT  0.185 1.955 0.445 2.455 ;
        END
        AntennaDiffArea 1.504 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.655 1.085 3.915 1.395 ;
        RECT  2.770 1.085 3.655 1.245 ;
        RECT  2.315 1.085 2.770 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.425 3.275 1.950 ;
        RECT  2.890 1.740 2.950 1.950 ;
        END
        AntennaGateArea 0.3952 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.170 1.005 1.495 1.395 ;
        RECT  0.855 0.920 1.170 1.395 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.200 2.070 1.775 ;
        RECT  0.615 1.615 1.700 1.775 ;
        RECT  0.355 1.220 0.615 1.775 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 -0.130 4.510 0.130 ;
        RECT  1.625 -0.130 1.885 0.400 ;
        RECT  0.000 -0.130 1.625 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.810 2.740 4.510 3.000 ;
        RECT  3.550 2.490 3.810 3.000 ;
        RECT  2.720 2.740 3.550 3.000 ;
        RECT  2.460 2.490 2.720 3.000 ;
        RECT  1.305 2.740 2.460 3.000 ;
        RECT  1.045 2.315 1.305 3.000 ;
        RECT  0.000 2.740 1.045 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.435 0.405 4.105 0.565 ;
        RECT  2.175 0.405 2.435 0.905 ;
        RECT  0.390 0.580 2.175 0.740 ;
        RECT  0.130 0.385 0.390 0.985 ;
    END
END OAI211X4MTH

MACRO OAI211X8MTH
    CLASS CORE ;
    FOREIGN OAI211X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.480 1.495 8.510 2.315 ;
        RECT  8.175 0.745 8.480 2.315 ;
        RECT  5.215 0.745 8.175 0.905 ;
        RECT  7.440 1.965 8.175 2.315 ;
        RECT  7.090 1.965 7.440 2.480 ;
        RECT  6.450 2.130 7.090 2.480 ;
        RECT  6.100 2.015 6.450 2.480 ;
        RECT  0.395 2.015 6.100 2.365 ;
        RECT  0.135 1.765 0.395 2.365 ;
        END
        AntennaDiffArea 3.002 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.835 1.085 7.995 1.405 ;
        RECT  6.475 1.085 7.835 1.245 ;
        RECT  5.875 1.085 6.475 1.345 ;
        RECT  4.820 1.085 5.875 1.245 ;
        RECT  4.415 1.085 4.820 1.580 ;
        END
        AntennaGateArea 0.7982 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.910 1.425 7.305 1.725 ;
        RECT  6.705 1.425 6.910 1.950 ;
        RECT  6.620 1.525 6.705 1.950 ;
        RECT  5.645 1.525 6.620 1.685 ;
        RECT  5.045 1.425 5.645 1.685 ;
        END
        AntennaGateArea 0.7904 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 0.985 3.440 1.435 ;
        RECT  1.515 0.985 3.180 1.145 ;
        RECT  1.130 0.985 1.515 1.445 ;
        RECT  0.915 0.880 1.130 1.445 ;
        END
        AntennaGateArea 0.8216 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.985 1.315 4.145 1.795 ;
        RECT  2.400 1.635 3.985 1.795 ;
        RECT  2.100 1.330 2.400 1.795 ;
        RECT  0.735 1.635 2.100 1.795 ;
        RECT  0.575 1.220 0.735 1.795 ;
        RECT  0.305 1.220 0.575 1.480 ;
        END
        AntennaGateArea 0.8216 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.475 -0.130 8.610 0.130 ;
        RECT  8.215 -0.130 8.475 0.300 ;
        RECT  2.985 -0.130 8.215 0.130 ;
        RECT  2.725 -0.130 2.985 0.465 ;
        RECT  0.935 -0.130 2.725 0.130 ;
        RECT  0.675 -0.130 0.935 0.360 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.935 2.740 8.610 3.000 ;
        RECT  7.675 2.495 7.935 3.000 ;
        RECT  5.865 2.740 7.675 3.000 ;
        RECT  5.605 2.545 5.865 3.000 ;
        RECT  3.225 2.740 5.605 3.000 ;
        RECT  2.965 2.545 3.225 3.000 ;
        RECT  1.280 2.740 2.965 3.000 ;
        RECT  1.020 2.545 1.280 3.000 ;
        RECT  0.000 2.740 1.020 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.590 0.405 7.965 0.565 ;
        RECT  4.330 0.405 4.590 0.905 ;
        RECT  1.485 0.645 4.330 0.805 ;
        RECT  1.325 0.540 1.485 0.805 ;
        RECT  0.385 0.540 1.325 0.700 ;
        RECT  0.125 0.410 0.385 1.010 ;
    END
END OAI211X8MTH

MACRO OAI211XLMTH
    CLASS CORE ;
    FOREIGN OAI211XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.905 0.785 2.295 0.945 ;
        RECT  1.905 1.740 1.990 1.950 ;
        RECT  1.745 0.785 1.905 1.950 ;
        RECT  1.700 1.740 1.745 1.950 ;
        RECT  0.125 1.790 1.700 1.950 ;
        END
        AntennaDiffArea 0.365 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.235 1.175 1.565 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 1.125 2.360 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 1.055 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.250 2.130 0.760 2.370 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.175 -0.130 2.460 0.130 ;
        RECT  1.575 -0.130 2.175 0.405 ;
        RECT  1.320 -0.130 1.575 0.130 ;
        RECT  0.720 -0.130 1.320 0.405 ;
        RECT  0.000 -0.130 0.720 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  2.075 2.110 2.335 3.000 ;
        RECT  1.790 2.740 2.075 3.000 ;
        RECT  1.530 2.570 1.790 3.000 ;
        RECT  1.245 2.740 1.530 3.000 ;
        RECT  0.985 2.130 1.245 3.000 ;
        RECT  0.000 2.740 0.985 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.125 0.735 1.405 0.995 ;
    END
END OAI211XLMTH

MACRO OAI21BX1MTH
    CLASS CORE ;
    FOREIGN OAI21BX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 0.935 1.855 1.095 ;
        RECT  1.560 0.935 1.635 1.550 ;
        RECT  1.475 0.935 1.560 2.235 ;
        RECT  1.330 1.290 1.475 2.235 ;
        RECT  0.985 1.975 1.330 2.235 ;
        END
        AntennaDiffArea 0.355 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.815 1.280 1.995 1.990 ;
        RECT  1.740 1.700 1.815 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.565 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.745 1.290 1.150 1.700 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.690 -0.130 2.460 0.130 ;
        RECT  0.750 -0.130 1.690 0.250 ;
        RECT  0.000 -0.130 0.750 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 2.740 2.460 3.000 ;
        RECT  1.525 2.415 1.785 3.000 ;
        RECT  0.385 2.740 1.525 3.000 ;
        RECT  0.125 1.830 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.175 0.310 2.335 2.380 ;
        RECT  2.075 0.310 2.175 0.670 ;
        RECT  2.120 2.120 2.175 2.380 ;
        RECT  1.255 0.510 2.075 0.670 ;
        RECT  1.135 0.850 1.295 1.110 ;
        RECT  0.390 0.850 1.135 1.010 ;
        RECT  0.130 0.735 0.390 1.010 ;
    END
END OAI21BX1MTH

MACRO OAI21BX2MTH
    CLASS CORE ;
    FOREIGN OAI21BX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.675 0.385 1.950 1.185 ;
        RECT  1.530 1.025 1.675 1.185 ;
        RECT  1.370 1.025 1.530 2.425 ;
        RECT  1.155 1.825 1.370 2.425 ;
        END
        AntennaDiffArea 0.585 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.215 2.705 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.635 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.840 1.160 1.190 1.645 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.785 -0.130 3.280 0.130 ;
        RECT  2.445 -0.130 2.785 0.300 ;
        RECT  2.185 -0.130 2.445 1.025 ;
        RECT  0.860 -0.130 2.185 0.130 ;
        RECT  0.600 -0.130 0.860 0.615 ;
        RECT  0.000 -0.130 0.600 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.650 2.740 3.280 3.000 ;
        RECT  1.970 2.440 2.650 3.000 ;
        RECT  1.710 2.100 1.970 3.000 ;
        RECT  0.550 2.740 1.710 3.000 ;
        RECT  0.290 1.760 0.550 3.000 ;
        RECT  0.000 2.740 0.290 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.900 0.765 3.060 1.920 ;
        RECT  2.735 0.765 2.900 1.025 ;
        RECT  1.970 1.760 2.900 1.920 ;
        RECT  1.710 1.365 1.970 1.920 ;
        RECT  1.200 0.550 1.425 0.810 ;
        RECT  1.040 0.550 1.200 0.960 ;
        RECT  0.385 0.800 1.040 0.960 ;
        RECT  0.125 0.360 0.385 0.960 ;
    END
END OAI21BX2MTH

MACRO OAI21BX4MTH
    CLASS CORE ;
    FOREIGN OAI21BX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.805 0.765 2.890 1.025 ;
        RECT  2.560 0.765 2.805 2.400 ;
        RECT  1.325 2.060 2.560 2.240 ;
        RECT  1.065 2.060 1.325 2.320 ;
        END
        AntennaDiffArea 0.948 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.410 1.220 4.000 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.220 2.105 1.880 ;
        RECT  0.675 1.720 1.700 1.880 ;
        RECT  0.515 1.220 0.675 1.880 ;
        RECT  0.415 1.220 0.515 1.480 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.220 1.495 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.825 -0.130 4.510 0.130 ;
        RECT  3.565 -0.130 3.825 0.515 ;
        RECT  1.860 -0.130 3.565 0.130 ;
        RECT  1.600 -0.130 1.860 0.700 ;
        RECT  0.000 -0.130 1.600 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.405 2.740 4.510 3.000 ;
        RECT  3.145 2.100 3.405 3.000 ;
        RECT  2.265 2.740 3.145 3.000 ;
        RECT  2.005 2.420 2.265 3.000 ;
        RECT  0.465 2.740 2.005 3.000 ;
        RECT  0.205 2.060 0.465 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.225 0.630 4.385 1.920 ;
        RECT  4.125 0.630 4.225 0.890 ;
        RECT  3.950 1.760 4.225 1.920 ;
        RECT  3.690 1.760 3.950 2.360 ;
        RECT  3.145 1.760 3.690 1.920 ;
        RECT  3.300 0.765 3.400 1.025 ;
        RECT  3.140 0.405 3.300 1.025 ;
        RECT  2.985 1.220 3.145 1.920 ;
        RECT  2.330 0.405 3.140 0.565 ;
        RECT  2.170 0.405 2.330 1.040 ;
        RECT  1.335 0.880 2.170 1.040 ;
        RECT  1.075 0.395 1.335 1.040 ;
        RECT  0.390 0.880 1.075 1.040 ;
        RECT  0.130 0.410 0.390 1.040 ;
    END
END OAI21BX4MTH

MACRO OAI21BX8MTH
    CLASS CORE ;
    FOREIGN OAI21BX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.915 0.785 6.105 1.135 ;
        RECT  5.845 1.725 6.105 2.330 ;
        RECT  5.025 1.725 5.845 2.075 ;
        RECT  4.915 1.725 5.025 2.255 ;
        RECT  4.565 0.785 4.915 2.255 ;
        RECT  3.625 1.905 4.565 2.255 ;
        RECT  3.365 1.905 3.625 2.515 ;
        RECT  1.565 1.905 3.365 2.255 ;
        RECT  1.305 1.905 1.565 2.505 ;
        END
        AntennaDiffArea 1.86 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.730 1.220 7.325 1.555 ;
        END
        AntennaGateArea 0.2054 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.015 1.265 4.275 1.685 ;
        RECT  2.810 1.525 4.015 1.685 ;
        RECT  2.135 1.260 2.810 1.685 ;
        RECT  0.725 1.525 2.135 1.685 ;
        RECT  0.465 1.220 0.725 1.685 ;
        END
        AntennaGateArea 0.8216 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.355 1.185 3.795 1.345 ;
        RECT  3.195 0.920 3.355 1.345 ;
        RECT  1.735 0.920 3.195 1.080 ;
        RECT  1.135 0.920 1.735 1.345 ;
        END
        AntennaGateArea 0.8216 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.125 -0.130 7.790 0.130 ;
        RECT  6.865 -0.130 7.125 1.025 ;
        RECT  3.025 -0.130 6.865 0.130 ;
        RECT  2.765 -0.130 3.025 0.400 ;
        RECT  0.935 -0.130 2.765 0.130 ;
        RECT  0.675 -0.130 0.935 0.400 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.055 2.740 7.790 3.000 ;
        RECT  6.455 2.110 7.055 3.000 ;
        RECT  5.565 2.740 6.455 3.000 ;
        RECT  5.305 2.255 5.565 3.000 ;
        RECT  4.485 2.740 5.305 3.000 ;
        RECT  4.225 2.480 4.485 3.000 ;
        RECT  2.765 2.740 4.225 3.000 ;
        RECT  2.165 2.480 2.765 3.000 ;
        RECT  0.735 2.740 2.165 3.000 ;
        RECT  0.135 1.915 0.735 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.505 0.385 7.665 2.400 ;
        RECT  7.405 0.385 7.505 0.985 ;
        RECT  7.405 1.735 7.505 2.400 ;
        RECT  6.465 1.735 7.405 1.895 ;
        RECT  6.355 0.405 6.615 1.005 ;
        RECT  6.305 1.345 6.465 1.895 ;
        RECT  4.315 0.405 6.355 0.565 ;
        RECT  5.165 1.345 6.305 1.505 ;
        RECT  4.155 0.405 4.315 0.740 ;
        RECT  3.575 0.580 4.155 0.740 ;
        RECT  3.315 0.450 3.575 0.740 ;
        RECT  2.475 0.580 3.315 0.740 ;
        RECT  2.215 0.450 2.475 0.740 ;
        RECT  1.485 0.580 2.215 0.740 ;
        RECT  1.225 0.445 1.485 0.740 ;
        RECT  0.385 0.580 1.225 0.740 ;
        RECT  0.125 0.385 0.385 0.985 ;
    END
END OAI21BX8MTH

MACRO OAI21BXLMTH
    CLASS CORE ;
    FOREIGN OAI21BXLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 0.935 1.885 1.095 ;
        RECT  1.540 0.935 1.665 1.525 ;
        RECT  1.505 0.935 1.540 2.090 ;
        RECT  1.330 1.365 1.505 2.090 ;
        RECT  0.985 1.830 1.330 2.090 ;
        END
        AntennaDiffArea 0.238 ;
    END Y
    PIN B0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 1.275 2.030 1.990 ;
        RECT  1.740 1.700 1.845 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END B0N
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.365 1.205 0.440 1.520 ;
        RECT  0.100 1.205 0.365 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.805 1.310 1.055 1.570 ;
        RECT  0.620 1.310 0.805 1.990 ;
        RECT  0.510 1.690 0.620 1.990 ;
        END
        AntennaGateArea 0.0858 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 -0.130 2.460 0.130 ;
        RECT  1.505 -0.130 1.765 0.330 ;
        RECT  1.065 -0.130 1.505 0.130 ;
        RECT  0.125 -0.130 1.065 0.415 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 2.740 2.460 3.000 ;
        RECT  0.810 2.450 1.750 3.000 ;
        RECT  0.385 2.740 0.810 3.000 ;
        RECT  0.125 2.120 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.210 0.310 2.370 2.380 ;
        RECT  2.075 0.310 2.210 0.670 ;
        RECT  2.060 2.170 2.210 2.380 ;
        RECT  1.255 0.510 2.075 0.670 ;
        RECT  1.165 0.850 1.325 1.145 ;
        RECT  0.385 0.850 1.165 1.010 ;
        RECT  0.125 0.740 0.385 1.010 ;
    END
END OAI21BXLMTH

MACRO OAI21X1MTH
    CLASS CORE ;
    FOREIGN OAI21X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.725 1.950 2.085 ;
        RECT  1.715 0.725 1.740 0.985 ;
        RECT  0.985 1.825 1.740 2.085 ;
        END
        AntennaDiffArea 0.358 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.115 1.560 1.645 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.165 0.615 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.115 1.130 1.625 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 -0.130 2.050 0.130 ;
        RECT  1.095 -0.130 1.695 0.415 ;
        RECT  0.810 -0.130 1.095 0.130 ;
        RECT  0.210 -0.130 0.810 0.415 ;
        RECT  0.000 -0.130 0.210 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 2.740 2.050 3.000 ;
        RECT  1.525 2.335 1.785 3.000 ;
        RECT  0.385 2.740 1.525 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.125 0.775 1.415 0.935 ;
    END
END OAI21X1MTH

MACRO OAI21X2MTH
    CLASS CORE ;
    FOREIGN OAI21X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.355 1.950 2.085 ;
        RECT  1.665 0.355 1.740 0.955 ;
        RECT  1.245 1.825 1.740 2.085 ;
        RECT  0.985 1.825 1.245 2.425 ;
        END
        AntennaDiffArea 0.571 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.135 1.555 1.645 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.165 0.615 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.795 1.135 1.130 1.625 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.895 -0.130 2.050 0.130 ;
        RECT  0.635 -0.130 0.895 0.565 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 2.740 2.050 3.000 ;
        RECT  1.525 2.335 1.785 3.000 ;
        RECT  0.385 2.740 1.525 3.000 ;
        RECT  0.125 1.835 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.155 0.355 1.415 0.955 ;
        RECT  0.385 0.795 1.155 0.955 ;
        RECT  0.125 0.355 0.385 0.955 ;
    END
END OAI21X2MTH

MACRO OAI21X3MTH
    CLASS CORE ;
    FOREIGN OAI21X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 1.290 3.180 1.920 ;
        RECT  2.965 0.815 3.125 1.920 ;
        RECT  2.765 0.815 2.965 0.975 ;
        RECT  2.905 1.760 2.965 1.920 ;
        RECT  2.645 1.760 2.905 2.360 ;
        RECT  1.185 2.045 2.645 2.305 ;
        END
        AntennaDiffArea 0.72 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.355 1.220 2.770 1.580 ;
        END
        AntennaGateArea 0.312 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.290 2.175 1.580 ;
        RECT  1.740 1.290 1.900 1.785 ;
        RECT  0.675 1.625 1.740 1.785 ;
        RECT  0.515 1.220 0.675 1.785 ;
        END
        AntennaGateArea 0.312 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.170 1.185 1.555 1.445 ;
        RECT  0.880 0.920 1.170 1.445 ;
        END
        AntennaGateArea 0.312 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 -0.130 3.690 0.130 ;
        RECT  1.735 -0.130 1.995 0.625 ;
        RECT  0.000 -0.130 1.735 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 2.740 3.690 3.000 ;
        RECT  3.185 2.100 3.445 3.000 ;
        RECT  2.335 2.740 3.185 3.000 ;
        RECT  2.075 2.495 2.335 3.000 ;
        RECT  0.575 2.740 2.075 3.000 ;
        RECT  0.315 2.030 0.575 3.000 ;
        RECT  0.000 2.740 0.315 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.305 0.475 3.565 0.830 ;
        RECT  2.545 0.475 3.305 0.635 ;
        RECT  2.285 0.475 2.545 0.975 ;
        RECT  1.510 0.815 2.285 0.975 ;
        RECT  1.350 0.580 1.510 0.975 ;
        RECT  0.385 0.580 1.350 0.740 ;
        RECT  0.125 0.580 0.385 0.910 ;
    END
END OAI21X3MTH

MACRO OAI21X4MTH
    CLASS CORE ;
    FOREIGN OAI21X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.150 1.290 3.210 1.945 ;
        RECT  2.970 0.805 3.150 1.945 ;
        RECT  2.795 0.805 2.970 0.985 ;
        RECT  2.945 1.765 2.970 1.945 ;
        RECT  2.685 1.765 2.945 2.420 ;
        RECT  1.175 2.060 2.685 2.320 ;
        END
        AntennaDiffArea 0.948 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.285 1.220 2.775 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 1.230 2.095 1.490 ;
        RECT  1.835 1.230 1.995 1.880 ;
        RECT  0.765 1.720 1.835 1.880 ;
        RECT  0.440 1.290 0.765 1.880 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.005 1.175 1.605 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 -0.130 3.690 0.130 ;
        RECT  1.725 -0.130 1.985 0.640 ;
        RECT  0.905 -0.130 1.725 0.130 ;
        RECT  0.645 -0.130 0.905 0.640 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.485 2.740 3.690 3.000 ;
        RECT  3.225 2.215 3.485 3.000 ;
        RECT  2.350 2.740 3.225 3.000 ;
        RECT  2.090 2.525 2.350 3.000 ;
        RECT  0.555 2.740 2.090 3.000 ;
        RECT  0.295 2.185 0.555 3.000 ;
        RECT  0.000 2.740 0.295 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.355 0.380 3.565 0.980 ;
        RECT  2.545 0.380 3.355 0.540 ;
        RECT  2.285 0.380 2.545 0.980 ;
        RECT  1.425 0.820 2.285 0.980 ;
        RECT  1.165 0.380 1.425 0.980 ;
        RECT  0.385 0.820 1.165 0.980 ;
        RECT  0.125 0.380 0.385 0.980 ;
    END
END OAI21X4MTH

MACRO OAI21X6MTH
    CLASS CORE ;
    FOREIGN OAI21X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 0.400 5.205 1.665 ;
        RECT  4.765 0.760 4.945 1.665 ;
        RECT  4.495 0.760 4.765 2.390 ;
        RECT  3.895 0.760 4.495 1.030 ;
        RECT  4.435 1.760 4.495 2.390 ;
        RECT  3.675 1.760 4.435 2.050 ;
        RECT  3.385 1.760 3.675 2.405 ;
        RECT  1.465 1.915 3.385 2.205 ;
        RECT  1.205 1.915 1.465 2.515 ;
        END
        AntennaDiffArea 1.529 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.755 1.220 4.305 1.580 ;
        END
        AntennaGateArea 0.6162 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.315 2.825 1.695 ;
        RECT  0.700 1.535 1.885 1.695 ;
        RECT  0.540 1.215 0.700 1.695 ;
        RECT  0.440 1.215 0.540 1.475 ;
        END
        AntennaGateArea 0.6162 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.285 0.920 3.445 1.575 ;
        RECT  1.635 0.920 3.285 1.080 ;
        RECT  0.880 0.920 1.635 1.355 ;
        END
        AntennaGateArea 0.6162 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.130 5.330 0.130 ;
        RECT  2.865 -0.130 3.125 0.385 ;
        RECT  2.025 -0.130 2.865 0.130 ;
        RECT  1.765 -0.130 2.025 0.390 ;
        RECT  0.000 -0.130 1.765 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 2.740 5.330 3.000 ;
        RECT  4.945 1.915 5.205 3.000 ;
        RECT  4.185 2.740 4.945 3.000 ;
        RECT  3.925 2.230 4.185 3.000 ;
        RECT  2.750 2.740 3.925 3.000 ;
        RECT  2.150 2.490 2.750 3.000 ;
        RECT  0.605 2.740 2.150 3.000 ;
        RECT  0.345 1.965 0.605 3.000 ;
        RECT  0.000 2.740 0.345 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.675 0.410 4.695 0.570 ;
        RECT  3.415 0.410 3.675 0.740 ;
        RECT  2.575 0.580 3.415 0.740 ;
        RECT  2.315 0.480 2.575 0.740 ;
        RECT  1.475 0.580 2.315 0.740 ;
        RECT  1.215 0.480 1.475 0.740 ;
        RECT  0.390 0.580 1.215 0.740 ;
        RECT  0.130 0.375 0.390 0.975 ;
    END
END OAI21X6MTH

MACRO OAI21X8MTH
    CLASS CORE ;
    FOREIGN OAI21X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.605 0.785 5.955 2.370 ;
        RECT  5.360 0.785 5.605 2.110 ;
        RECT  4.645 0.785 5.360 1.090 ;
        RECT  4.885 1.760 5.360 2.110 ;
        RECT  4.535 1.760 4.885 2.360 ;
        RECT  3.295 1.910 4.535 2.260 ;
        RECT  3.035 1.910 3.295 2.515 ;
        RECT  1.325 1.910 3.035 2.260 ;
        RECT  1.065 1.910 1.325 2.515 ;
        END
        AntennaDiffArea 1.956 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 1.270 5.160 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.745 1.315 4.005 1.690 ;
        RECT  2.500 1.530 3.745 1.690 ;
        RECT  1.885 1.315 2.500 1.690 ;
        RECT  0.675 1.530 1.885 1.690 ;
        RECT  0.415 1.220 0.675 1.690 ;
        END
        AntennaGateArea 0.8216 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 1.185 3.415 1.345 ;
        RECT  2.750 0.975 2.910 1.345 ;
        RECT  1.495 0.975 2.750 1.135 ;
        RECT  1.170 0.975 1.495 1.345 ;
        RECT  0.880 0.920 1.170 1.345 ;
        END
        AntennaGateArea 0.8216 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.865 -0.130 6.560 0.130 ;
        RECT  3.605 -0.130 3.865 0.565 ;
        RECT  1.865 -0.130 3.605 0.130 ;
        RECT  1.605 -0.130 1.865 0.400 ;
        RECT  0.000 -0.130 1.605 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.405 2.740 6.560 3.000 ;
        RECT  6.145 1.890 6.405 3.000 ;
        RECT  5.355 2.740 6.145 3.000 ;
        RECT  5.095 2.295 5.355 3.000 ;
        RECT  4.280 2.740 5.095 3.000 ;
        RECT  4.020 2.505 4.280 3.000 ;
        RECT  2.290 2.740 4.020 3.000 ;
        RECT  2.030 2.505 2.290 3.000 ;
        RECT  0.465 2.740 2.030 3.000 ;
        RECT  0.205 1.915 0.465 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.175 0.405 6.435 1.005 ;
        RECT  4.395 0.405 6.175 0.565 ;
        RECT  4.135 0.355 4.395 0.955 ;
        RECT  3.355 0.795 4.135 0.955 ;
        RECT  3.095 0.345 3.355 0.955 ;
        RECT  2.415 0.345 3.095 0.505 ;
        RECT  2.155 0.345 2.415 0.740 ;
        RECT  0.390 0.580 2.155 0.740 ;
        RECT  0.130 0.370 0.390 0.970 ;
    END
END OAI21X8MTH

MACRO OAI21XLMTH
    CLASS CORE ;
    FOREIGN OAI21XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.900 1.700 1.950 1.990 ;
        RECT  1.740 0.335 1.900 1.990 ;
        RECT  1.640 0.335 1.740 0.595 ;
        RECT  1.015 1.760 1.740 1.920 ;
        END
        AntennaDiffArea 0.363 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.205 1.205 1.560 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.330 1.205 0.355 1.580 ;
        RECT  0.100 1.205 0.330 1.840 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.865 1.205 1.025 1.465 ;
        RECT  0.720 1.305 0.865 1.465 ;
        RECT  0.560 1.305 0.720 1.990 ;
        RECT  0.510 1.700 0.560 1.990 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 -0.130 2.050 0.130 ;
        RECT  0.335 -0.130 1.275 0.515 ;
        RECT  0.000 -0.130 0.335 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.845 2.740 2.050 3.000 ;
        RECT  1.585 2.180 1.845 3.000 ;
        RECT  1.295 2.740 1.585 3.000 ;
        RECT  0.695 2.390 1.295 3.000 ;
        RECT  0.385 2.740 0.695 3.000 ;
        RECT  0.125 2.180 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.175 0.765 1.435 1.025 ;
        RECT  0.385 0.865 1.175 1.025 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END OAI21XLMTH

MACRO OAI221X1MTH
    CLASS CORE ;
    FOREIGN OAI221X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.005 0.705 3.180 2.035 ;
        RECT  2.895 0.705 3.005 0.965 ;
        RECT  2.970 1.700 3.005 2.035 ;
        RECT  0.490 1.875 2.970 2.035 ;
        RECT  0.230 1.875 0.490 2.135 ;
        END
        AntennaDiffArea 0.605 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.790 1.140 2.825 1.480 ;
        RECT  2.540 1.140 2.790 1.695 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.810 1.220 1.150 1.690 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.220 0.630 1.590 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.180 1.875 1.685 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 1.175 2.360 1.690 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 -0.130 3.280 0.130 ;
        RECT  2.865 -0.130 3.125 0.330 ;
        RECT  1.175 -0.130 2.865 0.130 ;
        RECT  0.235 -0.130 1.175 0.410 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.125 2.740 3.280 3.000 ;
        RECT  2.865 2.215 3.125 3.000 ;
        RECT  1.505 2.740 2.865 3.000 ;
        RECT  1.245 2.215 1.505 3.000 ;
        RECT  0.000 2.740 1.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.580 0.735 2.215 0.995 ;
    END
END OAI221X1MTH

MACRO OAI221X2MTH
    CLASS CORE ;
    FOREIGN OAI221X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 0.385 3.590 1.920 ;
        RECT  3.285 0.385 3.345 0.985 ;
        RECT  2.515 1.760 3.345 1.920 ;
        RECT  2.255 1.760 2.515 2.360 ;
        RECT  0.550 1.925 2.255 2.085 ;
        RECT  0.290 1.820 0.550 2.420 ;
        END
        AntennaDiffArea 0.867 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.220 3.145 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 1.165 1.150 1.735 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.320 1.160 0.720 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.160 1.775 1.725 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 1.135 2.380 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.935 -0.130 3.690 0.130 ;
        RECT  0.675 -0.130 0.935 0.640 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.395 2.740 3.690 3.000 ;
        RECT  2.795 2.100 3.395 3.000 ;
        RECT  1.530 2.740 2.795 3.000 ;
        RECT  1.270 2.280 1.530 3.000 ;
        RECT  0.000 2.740 1.270 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.775 0.355 3.035 0.955 ;
        RECT  1.745 0.795 2.775 0.955 ;
        RECT  2.265 0.355 2.525 0.615 ;
        RECT  1.485 0.455 2.265 0.615 ;
        RECT  1.225 0.455 1.485 0.980 ;
        RECT  0.385 0.820 1.225 0.980 ;
        RECT  0.125 0.375 0.385 0.980 ;
    END
END OAI221X2MTH

MACRO OAI221X4MTH
    CLASS CORE ;
    FOREIGN OAI221X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.805 0.805 6.050 2.405 ;
        RECT  5.240 0.805 5.805 0.985 ;
        RECT  5.765 1.720 5.805 2.405 ;
        RECT  4.565 1.720 5.765 1.900 ;
        RECT  4.305 1.720 4.565 2.405 ;
        RECT  2.380 2.130 4.305 2.310 ;
        RECT  2.120 1.925 2.380 2.475 ;
        RECT  0.505 1.925 2.120 2.105 ;
        RECT  0.245 1.925 0.505 2.460 ;
        END
        AntennaDiffArea 1.688 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.645 1.220 5.585 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 0.920 1.495 1.405 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.220 2.135 1.745 ;
        RECT  0.675 1.585 1.700 1.745 ;
        RECT  0.415 1.220 0.675 1.745 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.210 3.685 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.090 1.220 4.345 1.480 ;
        RECT  3.930 1.220 4.090 1.880 ;
        RECT  2.770 1.720 3.930 1.880 ;
        RECT  2.560 1.220 2.770 1.880 ;
        RECT  2.355 1.220 2.560 1.480 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 -0.130 6.150 0.130 ;
        RECT  1.625 -0.130 1.885 0.400 ;
        RECT  0.000 -0.130 1.625 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.470 2.740 6.150 3.000 ;
        RECT  4.870 2.145 5.470 3.000 ;
        RECT  3.655 2.740 4.870 3.000 ;
        RECT  3.055 2.490 3.655 3.000 ;
        RECT  1.405 2.740 3.055 3.000 ;
        RECT  1.145 2.290 1.405 3.000 ;
        RECT  0.000 2.740 1.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.765 0.365 6.025 0.625 ;
        RECT  5.005 0.465 5.765 0.625 ;
        RECT  4.845 0.465 5.005 1.025 ;
        RECT  4.745 0.745 4.845 1.025 ;
        RECT  2.695 0.745 4.745 0.905 ;
        RECT  2.435 0.405 4.525 0.565 ;
        RECT  2.175 0.405 2.435 0.905 ;
        RECT  1.335 0.580 2.175 0.740 ;
        RECT  1.075 0.480 1.335 0.740 ;
        RECT  0.390 0.580 1.075 0.740 ;
        RECT  0.130 0.385 0.390 0.985 ;
    END
END OAI221X4MTH

MACRO OAI221XLMTH
    CLASS CORE ;
    FOREIGN OAI221XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 0.325 3.180 1.920 ;
        RECT  2.895 0.325 2.970 0.585 ;
        RECT  0.190 1.760 2.970 1.920 ;
        END
        AntennaDiffArea 0.492 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 2.100 2.665 2.400 ;
        END
        AntennaGateArea 0.0702 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.810 1.220 1.150 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.220 0.620 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.220 1.875 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.095 1.220 2.770 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.155 -0.130 3.280 0.130 ;
        RECT  0.215 -0.130 1.155 0.515 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.105 2.740 3.280 3.000 ;
        RECT  2.845 2.170 3.105 3.000 ;
        RECT  2.570 2.740 2.845 3.000 ;
        RECT  1.630 2.620 2.570 3.000 ;
        RECT  1.320 2.740 1.630 3.000 ;
        RECT  1.060 2.100 1.320 3.000 ;
        RECT  0.680 2.740 1.060 3.000 ;
        RECT  0.420 2.620 0.680 3.000 ;
        RECT  0.000 2.740 0.420 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.565 0.765 2.215 1.025 ;
    END
END OAI221XLMTH

MACRO OAI222X1MTH
    CLASS CORE ;
    FOREIGN OAI222X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 1.700 3.180 2.290 ;
        RECT  2.970 0.735 3.155 2.290 ;
        RECT  2.900 0.735 2.970 0.995 ;
        RECT  0.495 2.130 2.970 2.290 ;
        RECT  0.235 1.920 0.495 2.290 ;
        END
        AntennaDiffArea 0.669 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.335 1.010 3.600 1.605 ;
        END
        AntennaGateArea 0.1274 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 1.235 2.790 1.795 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 1.740 1.210 1.950 ;
        RECT  0.880 1.265 1.150 1.950 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.265 0.665 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.615 1.175 1.885 1.520 ;
        RECT  1.330 1.175 1.615 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 1.400 2.315 1.950 ;
        RECT  1.700 1.740 2.120 1.950 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.185 -0.130 3.690 0.130 ;
        RECT  0.245 -0.130 1.185 0.405 ;
        RECT  0.000 -0.130 0.245 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 2.740 3.690 3.000 ;
        RECT  3.255 2.455 3.515 3.000 ;
        RECT  1.505 2.740 3.255 3.000 ;
        RECT  1.245 2.470 1.505 3.000 ;
        RECT  0.000 2.740 1.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.585 0.735 2.225 0.995 ;
    END
END OAI222X1MTH

MACRO OAI222X2MTH
    CLASS CORE ;
    FOREIGN OAI222X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.745 4.000 2.005 ;
        RECT  3.205 0.745 3.790 0.905 ;
        RECT  2.830 1.845 3.790 2.005 ;
        RECT  2.330 1.845 2.830 2.445 ;
        RECT  0.395 1.845 2.330 2.005 ;
        RECT  0.135 1.845 0.395 2.445 ;
        END
        AntennaDiffArea 1.332 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.360 1.085 3.610 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.725 1.155 3.180 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.785 1.140 1.150 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.145 0.605 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.175 1.825 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.005 1.155 2.530 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.905 -0.130 4.100 0.130 ;
        RECT  0.645 -0.130 0.905 0.615 ;
        RECT  0.000 -0.130 0.645 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.815 2.740 4.100 3.000 ;
        RECT  3.555 2.185 3.815 3.000 ;
        RECT  1.595 2.740 3.555 3.000 ;
        RECT  0.995 2.185 1.595 3.000 ;
        RECT  0.000 2.740 0.995 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.955 0.405 3.975 0.565 ;
        RECT  2.795 0.405 2.955 0.975 ;
        RECT  1.945 0.815 2.795 0.975 ;
        RECT  2.205 0.375 2.465 0.565 ;
        RECT  1.425 0.375 2.205 0.535 ;
        RECT  1.685 0.715 1.945 0.975 ;
        RECT  1.165 0.375 1.425 0.955 ;
        RECT  0.385 0.795 1.165 0.955 ;
        RECT  0.125 0.355 0.385 0.955 ;
    END
END OAI222X2MTH

MACRO OAI222X4MTH
    CLASS CORE ;
    FOREIGN OAI222X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.070 0.745 7.280 1.990 ;
        RECT  5.425 0.745 7.070 0.905 ;
        RECT  6.865 1.810 7.070 1.990 ;
        RECT  6.635 1.810 6.865 2.415 ;
        RECT  4.915 2.130 6.635 2.310 ;
        RECT  4.315 1.880 4.915 2.480 ;
        RECT  2.530 2.130 4.315 2.310 ;
        RECT  2.270 1.965 2.530 2.465 ;
        RECT  0.655 1.965 2.270 2.145 ;
        RECT  0.395 1.965 0.655 2.465 ;
        END
        AntennaDiffArea 2.454 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.565 1.180 6.115 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.615 1.235 6.875 1.565 ;
        RECT  6.455 1.405 6.615 1.565 ;
        RECT  6.295 1.405 6.455 1.890 ;
        RECT  5.365 1.730 6.295 1.890 ;
        RECT  5.205 1.160 5.365 1.890 ;
        RECT  4.900 1.160 5.205 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 0.920 1.705 1.445 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 1.265 2.360 1.785 ;
        RECT  0.780 1.625 1.985 1.785 ;
        RECT  0.520 1.220 0.780 1.785 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.185 1.120 3.785 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.125 1.200 4.305 1.510 ;
        RECT  3.965 1.200 4.125 1.880 ;
        RECT  2.915 1.720 3.965 1.880 ;
        RECT  2.755 1.200 2.915 1.880 ;
        RECT  2.560 1.200 2.755 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.035 -0.130 7.380 0.130 ;
        RECT  1.775 -0.130 2.035 0.400 ;
        RECT  0.935 -0.130 1.775 0.130 ;
        RECT  0.675 -0.130 0.935 0.400 ;
        RECT  0.000 -0.130 0.675 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.915 2.740 7.380 3.000 ;
        RECT  5.655 2.490 5.915 3.000 ;
        RECT  3.550 2.740 5.655 3.000 ;
        RECT  3.290 2.490 3.550 3.000 ;
        RECT  1.535 2.740 3.290 3.000 ;
        RECT  1.275 2.335 1.535 3.000 ;
        RECT  0.000 2.740 1.275 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.175 0.405 7.215 0.565 ;
        RECT  4.915 0.405 5.175 0.905 ;
        RECT  2.845 0.745 4.915 0.905 ;
        RECT  2.585 0.405 4.665 0.565 ;
        RECT  2.325 0.405 2.585 0.740 ;
        RECT  1.485 0.580 2.325 0.740 ;
        RECT  1.225 0.480 1.485 0.740 ;
        RECT  0.390 0.580 1.225 0.740 ;
        RECT  0.130 0.385 0.390 0.985 ;
    END
END OAI222X4MTH

MACRO OAI222XLMTH
    CLASS CORE ;
    FOREIGN OAI222XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 1.700 3.180 2.290 ;
        RECT  2.970 0.765 3.155 2.290 ;
        RECT  2.910 0.765 2.970 1.025 ;
        RECT  0.495 2.130 2.970 2.290 ;
        RECT  0.235 1.770 0.495 2.290 ;
        END
        AntennaDiffArea 0.568 ;
    END Y
    PIN C1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.335 1.010 3.600 1.605 ;
        END
        AntennaGateArea 0.0858 ;
    END C1
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.505 1.235 2.790 1.725 ;
        END
        AntennaGateArea 0.0858 ;
    END C0
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.265 1.150 1.845 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.265 0.665 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.175 1.785 1.520 ;
        RECT  1.330 1.175 1.540 1.655 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.025 1.400 2.315 1.950 ;
        RECT  1.700 1.740 2.025 1.950 ;
        END
        AntennaGateArea 0.0858 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.165 -0.130 3.690 0.130 ;
        RECT  0.225 -0.130 1.165 0.405 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.515 2.740 3.690 3.000 ;
        RECT  2.915 2.505 3.515 3.000 ;
        RECT  1.565 2.740 2.915 3.000 ;
        RECT  0.625 2.480 1.565 3.000 ;
        RECT  0.000 2.740 0.625 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.955 0.735 2.215 1.025 ;
        RECT  0.825 0.735 1.955 0.895 ;
        RECT  0.565 0.735 0.825 1.025 ;
    END
END OAI222XLMTH

MACRO OAI22X1MTH
    CLASS CORE ;
    FOREIGN OAI22X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.970 1.350 2.130 ;
        RECT  0.970 1.290 1.130 2.130 ;
        RECT  0.915 1.290 0.970 1.580 ;
        RECT  0.855 1.290 0.915 1.450 ;
        RECT  0.695 0.760 0.855 1.450 ;
        RECT  0.525 0.760 0.695 1.020 ;
        END
        AntennaDiffArea 0.36 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.165 2.360 1.580 ;
        RECT  1.740 1.165 2.150 1.425 ;
        END
        AntennaGateArea 0.1235 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.630 1.950 1.990 ;
        RECT  1.520 1.630 1.740 1.790 ;
        RECT  1.310 1.280 1.520 1.790 ;
        END
        AntennaGateArea 0.1235 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.245 0.495 1.505 ;
        RECT  0.100 0.880 0.335 1.505 ;
        END
        AntennaGateArea 0.1235 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 2.395 1.180 2.555 ;
        RECT  0.565 1.700 0.725 2.555 ;
        RECT  0.510 1.700 0.565 1.990 ;
        END
        AntennaGateArea 0.1235 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.185 -0.130 2.460 0.130 ;
        RECT  1.585 -0.130 2.185 0.415 ;
        RECT  0.000 -0.130 1.585 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 2.740 2.460 3.000 ;
        RECT  1.950 2.170 2.210 3.000 ;
        RECT  0.385 2.740 1.950 3.000 ;
        RECT  0.125 2.180 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.075 0.725 2.335 0.985 ;
        RECT  1.295 0.825 2.075 0.985 ;
        RECT  1.035 0.725 1.295 0.985 ;
    END
END OAI22X1MTH

MACRO OAI22X2MTH
    CLASS CORE ;
    FOREIGN OAI22X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.155 1.840 1.540 2.440 ;
        RECT  0.695 1.840 1.155 2.000 ;
        RECT  0.695 0.815 0.895 0.975 ;
        RECT  0.535 0.815 0.695 2.000 ;
        END
        AntennaDiffArea 0.722 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 1.245 2.770 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.445 1.240 1.950 1.650 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.355 1.535 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.160 1.265 1.645 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.955 -0.130 2.870 0.130 ;
        RECT  1.695 -0.130 1.955 0.640 ;
        RECT  0.000 -0.130 1.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.730 2.740 2.870 3.000 ;
        RECT  2.130 1.760 2.730 3.000 ;
        RECT  0.485 2.740 2.130 3.000 ;
        RECT  0.225 2.180 0.485 3.000 ;
        RECT  0.000 2.740 0.225 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.245 0.380 2.505 0.980 ;
        RECT  1.405 0.820 2.245 0.980 ;
        RECT  1.145 0.380 1.405 0.980 ;
        RECT  0.385 0.380 1.145 0.540 ;
        RECT  0.125 0.380 0.385 0.680 ;
    END
END OAI22X2MTH

MACRO OAI22X4MTH
    CLASS CORE ;
    FOREIGN OAI22X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 1.700 4.545 2.360 ;
        RECT  2.360 2.060 4.200 2.240 ;
        RECT  2.200 1.830 2.360 2.430 ;
        RECT  0.535 2.060 2.200 2.240 ;
        RECT  0.330 0.795 1.915 0.975 ;
        RECT  0.330 1.915 0.535 2.515 ;
        RECT  0.150 0.795 0.330 2.515 ;
        END
        AntennaDiffArea 1.584 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.930 1.205 3.570 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.235 4.375 1.460 ;
        RECT  3.790 1.235 4.000 1.880 ;
        RECT  2.700 1.720 3.790 1.880 ;
        RECT  2.540 1.245 2.700 1.880 ;
        RECT  2.395 1.245 2.540 1.505 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.055 1.205 1.655 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 1.245 2.175 1.505 ;
        RECT  1.835 1.245 1.995 1.880 ;
        RECT  0.875 1.720 1.835 1.880 ;
        RECT  0.715 1.235 0.875 1.880 ;
        RECT  0.510 1.235 0.715 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.075 -0.130 4.920 0.130 ;
        RECT  3.815 -0.130 4.075 0.605 ;
        RECT  2.975 -0.130 3.815 0.130 ;
        RECT  2.715 -0.130 2.975 0.605 ;
        RECT  0.000 -0.130 2.715 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.685 2.740 4.920 3.000 ;
        RECT  3.085 2.460 3.685 3.000 ;
        RECT  1.465 2.740 3.085 3.000 ;
        RECT  1.205 2.460 1.465 3.000 ;
        RECT  0.000 2.740 1.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.365 0.355 4.625 0.955 ;
        RECT  3.525 0.795 4.365 0.955 ;
        RECT  3.265 0.355 3.525 0.955 ;
        RECT  2.425 0.795 3.265 0.955 ;
        RECT  2.165 0.355 2.425 0.955 ;
        RECT  0.125 0.455 2.165 0.615 ;
    END
END OAI22X4MTH

MACRO OAI22X8MTH
    CLASS CORE ;
    FOREIGN OAI22X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.480 1.085 8.510 1.785 ;
        RECT  8.245 0.745 8.480 2.505 ;
        RECT  4.655 0.745 8.245 0.905 ;
        RECT  8.025 1.905 8.245 2.505 ;
        RECT  6.975 1.905 8.025 2.255 ;
        RECT  6.685 1.905 6.975 2.520 ;
        RECT  6.030 2.170 6.685 2.520 ;
        RECT  5.675 2.015 6.030 2.520 ;
        RECT  4.350 2.015 5.675 2.365 ;
        RECT  4.090 1.765 4.350 2.365 ;
        RECT  0.425 2.015 4.090 2.365 ;
        RECT  0.165 1.965 0.425 2.465 ;
        END
        AntennaDiffArea 2.767 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.995 1.115 3.435 1.375 ;
        RECT  2.835 0.920 2.995 1.375 ;
        RECT  1.755 0.920 2.835 1.080 ;
        RECT  0.815 0.920 1.755 1.395 ;
        END
        AntennaGateArea 0.8216 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.780 1.235 4.065 1.495 ;
        RECT  3.620 1.235 3.780 1.735 ;
        RECT  2.595 1.575 3.620 1.735 ;
        RECT  1.995 1.315 2.595 1.735 ;
        RECT  0.595 1.575 1.995 1.735 ;
        RECT  0.435 1.220 0.595 1.735 ;
        RECT  0.335 1.220 0.435 1.480 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.960 1.425 7.560 1.685 ;
        RECT  6.500 1.525 6.960 1.685 ;
        RECT  6.210 1.525 6.500 1.950 ;
        RECT  5.600 1.525 6.210 1.685 ;
        RECT  5.000 1.425 5.600 1.685 ;
        END
        AntennaGateArea 0.7904 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.835 1.085 8.065 1.480 ;
        RECT  6.615 1.085 7.835 1.245 ;
        RECT  6.015 1.085 6.615 1.345 ;
        RECT  4.820 1.085 6.015 1.245 ;
        RECT  4.585 1.085 4.820 1.580 ;
        RECT  4.335 1.235 4.585 1.580 ;
        END
        AntennaGateArea 0.7904 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 -0.130 8.610 0.130 ;
        RECT  1.625 -0.130 1.885 0.400 ;
        RECT  0.000 -0.130 1.625 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.415 2.740 8.610 3.000 ;
        RECT  7.155 2.440 7.415 3.000 ;
        RECT  5.435 2.740 7.155 3.000 ;
        RECT  5.175 2.545 5.435 3.000 ;
        RECT  3.330 2.740 5.175 3.000 ;
        RECT  3.070 2.550 3.330 3.000 ;
        RECT  1.595 2.740 3.070 3.000 ;
        RECT  0.995 2.545 1.595 3.000 ;
        RECT  0.000 2.740 0.995 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.405 0.405 8.485 0.565 ;
        RECT  4.145 0.370 4.405 0.970 ;
        RECT  3.415 0.580 4.145 0.740 ;
        RECT  3.155 0.480 3.415 0.740 ;
        RECT  2.435 0.580 3.155 0.740 ;
        RECT  2.175 0.480 2.435 0.740 ;
        RECT  1.335 0.580 2.175 0.740 ;
        RECT  1.075 0.480 1.335 0.740 ;
        RECT  0.390 0.580 1.075 0.740 ;
        RECT  0.130 0.410 0.390 1.010 ;
    END
END OAI22X8MTH

MACRO OAI22XLMTH
    CLASS CORE ;
    FOREIGN OAI22XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.865 1.320 2.025 ;
        RECT  0.915 1.210 1.130 2.025 ;
        RECT  0.785 1.210 0.915 1.370 ;
        RECT  0.785 0.765 0.815 1.025 ;
        RECT  0.625 0.765 0.785 1.370 ;
        RECT  0.555 0.765 0.625 1.025 ;
        END
        AntennaDiffArea 0.296 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.185 2.360 1.580 ;
        RECT  1.740 1.185 2.150 1.345 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.525 1.950 1.990 ;
        RECT  1.520 1.525 1.740 1.685 ;
        RECT  1.310 1.215 1.520 1.685 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.335 1.260 0.445 1.520 ;
        RECT  0.100 0.880 0.335 1.520 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 2.235 1.120 2.395 ;
        RECT  0.565 1.700 0.725 2.395 ;
        RECT  0.510 1.700 0.565 1.990 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.185 -0.130 2.460 0.130 ;
        RECT  1.585 -0.130 2.185 0.515 ;
        RECT  0.000 -0.130 1.585 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 2.740 2.460 3.000 ;
        RECT  1.950 2.170 2.210 3.000 ;
        RECT  1.660 2.740 1.950 3.000 ;
        RECT  0.720 2.605 1.660 3.000 ;
        RECT  0.385 2.740 0.720 3.000 ;
        RECT  0.125 2.180 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.325 0.815 2.335 0.975 ;
        RECT  1.165 0.335 1.325 0.975 ;
        RECT  1.065 0.335 1.165 0.595 ;
    END
END OAI22XLMTH

MACRO OAI2B11X1MTH
    CLASS CORE ;
    FOREIGN OAI2B11X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 0.815 2.745 2.110 ;
        RECT  2.065 0.815 2.585 0.975 ;
        RECT  1.990 1.850 2.585 2.110 ;
        RECT  1.455 1.740 1.990 2.110 ;
        END
        AntennaDiffArea 0.577 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.145 3.180 1.665 ;
        END
        AntennaGateArea 0.1274 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.945 1.230 2.405 1.540 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.075 0.585 2.400 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.220 1.755 1.540 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.720 -0.130 3.280 0.130 ;
        RECT  0.780 -0.130 1.720 0.295 ;
        RECT  0.000 -0.130 0.780 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.130 2.740 3.280 3.000 ;
        RECT  2.940 1.850 3.130 3.000 ;
        RECT  2.755 2.740 2.940 3.000 ;
        RECT  1.815 2.555 2.755 3.000 ;
        RECT  1.635 2.740 1.815 3.000 ;
        RECT  0.695 2.555 1.635 3.000 ;
        RECT  0.000 2.740 0.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.940 0.475 3.100 0.965 ;
        RECT  1.385 0.475 2.940 0.635 ;
        RECT  1.225 0.475 1.385 0.995 ;
        RECT  1.125 0.735 1.225 0.995 ;
        RECT  0.805 1.230 1.065 1.490 ;
        RECT  0.385 1.330 0.805 1.490 ;
        RECT  0.225 0.765 0.385 1.895 ;
        RECT  0.125 0.765 0.225 1.025 ;
        RECT  0.125 1.735 0.225 1.895 ;
    END
END OAI2B11X1MTH

MACRO OAI2B11X2MTH
    CLASS CORE ;
    FOREIGN OAI2B11X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 1.700 2.770 1.990 ;
        RECT  2.635 0.770 2.720 1.990 ;
        RECT  2.560 0.770 2.635 2.430 ;
        RECT  2.065 0.770 2.560 0.930 ;
        RECT  2.375 1.770 2.560 2.430 ;
        RECT  1.725 1.770 2.375 1.930 ;
        RECT  1.465 1.770 1.725 2.030 ;
        END
        AntennaDiffArea 0.775 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.955 1.135 3.180 1.695 ;
        RECT  2.900 1.135 2.955 1.565 ;
        END
        AntennaGateArea 0.2054 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 1.225 2.380 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.110 0.605 2.405 ;
        END
        AntennaGateArea 0.0871 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.220 1.780 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 -0.130 3.280 0.130 ;
        RECT  1.665 -0.130 1.925 0.250 ;
        RECT  0.825 -0.130 1.665 0.130 ;
        RECT  0.225 -0.130 0.825 0.465 ;
        RECT  0.000 -0.130 0.225 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.145 2.740 3.280 3.000 ;
        RECT  2.885 2.145 3.145 3.000 ;
        RECT  2.125 2.740 2.885 3.000 ;
        RECT  1.865 2.255 2.125 3.000 ;
        RECT  0.850 2.740 1.865 3.000 ;
        RECT  0.250 2.585 0.850 3.000 ;
        RECT  0.000 2.740 0.250 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.905 0.350 3.150 0.955 ;
        RECT  1.375 0.430 2.905 0.590 ;
        RECT  1.115 0.380 1.375 0.980 ;
        RECT  0.800 1.225 1.060 1.485 ;
        RECT  0.385 1.325 0.800 1.485 ;
        RECT  0.225 0.765 0.385 1.925 ;
        RECT  0.125 0.765 0.225 1.025 ;
        RECT  0.125 1.705 0.225 1.925 ;
    END
END OAI2B11X2MTH

MACRO OAI2B11X4MTH
    CLASS CORE ;
    FOREIGN OAI2B11X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.060 0.770 5.240 2.280 ;
        RECT  4.020 0.770 5.060 0.950 ;
        RECT  5.020 1.700 5.060 2.280 ;
        RECT  4.655 2.100 5.020 2.280 ;
        RECT  4.395 2.100 4.655 2.360 ;
        RECT  3.655 2.100 4.395 2.280 ;
        RECT  3.395 2.100 3.655 2.360 ;
        RECT  1.865 2.100 3.395 2.280 ;
        RECT  1.605 2.100 1.865 2.360 ;
        END
        AntennaDiffArea 1.292 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.225 4.880 1.485 ;
        RECT  4.610 1.225 4.820 1.880 ;
        RECT  3.475 1.720 4.610 1.880 ;
        RECT  3.315 1.225 3.475 1.880 ;
        RECT  3.215 1.225 3.315 1.485 ;
        END
        AntennaGateArea 0.4108 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.750 1.225 4.250 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.620 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.225 2.075 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.050 -0.130 5.330 0.130 ;
        RECT  2.790 -0.130 3.050 0.515 ;
        RECT  0.925 -0.130 2.790 0.130 ;
        RECT  0.665 -0.130 0.925 0.685 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.205 2.740 5.330 3.000 ;
        RECT  4.945 2.460 5.205 3.000 ;
        RECT  3.090 2.740 4.945 3.000 ;
        RECT  2.490 2.480 3.090 3.000 ;
        RECT  0.990 2.740 2.490 3.000 ;
        RECT  0.730 2.100 0.990 3.000 ;
        RECT  0.000 2.740 0.730 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.450 0.430 5.110 0.590 ;
        RECT  3.230 0.430 3.450 0.965 ;
        RECT  2.500 0.805 3.230 0.965 ;
        RECT  2.580 1.225 2.680 1.485 ;
        RECT  2.420 1.225 2.580 1.920 ;
        RECT  2.240 0.365 2.500 0.965 ;
        RECT  1.150 1.760 2.420 1.920 ;
        RECT  1.475 0.805 2.240 0.965 ;
        RECT  1.215 0.365 1.475 0.965 ;
        RECT  1.035 1.225 1.150 1.920 ;
        RECT  0.875 0.865 1.035 1.920 ;
        RECT  0.385 0.865 0.875 1.025 ;
        RECT  0.450 1.760 0.875 1.920 ;
        RECT  0.190 1.760 0.450 2.360 ;
        RECT  0.125 0.605 0.385 1.025 ;
    END
END OAI2B11X4MTH

MACRO OAI2B11XLMTH
    CLASS CORE ;
    FOREIGN OAI2B11XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.580 0.815 2.740 1.980 ;
        RECT  2.085 0.815 2.580 0.975 ;
        RECT  1.455 1.720 2.580 1.980 ;
        END
        AntennaDiffArea 0.362 ;
    END Y
    PIN C0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.920 1.145 3.180 1.665 ;
        END
        AntennaGateArea 0.0702 ;
    END C0
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.945 1.225 2.400 1.540 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 2.100 0.585 2.400 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.220 1.755 1.540 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.340 -0.130 3.280 0.130 ;
        RECT  1.400 -0.130 2.340 0.295 ;
        RECT  1.140 -0.130 1.400 0.130 ;
        RECT  0.200 -0.130 1.140 0.295 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 2.740 3.280 3.000 ;
        RECT  2.035 2.570 2.975 3.000 ;
        RECT  1.815 2.740 2.035 3.000 ;
        RECT  0.875 2.570 1.815 3.000 ;
        RECT  0.000 2.740 0.875 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.895 0.335 3.155 0.635 ;
        RECT  1.345 0.475 2.895 0.635 ;
        RECT  1.185 0.475 1.345 0.940 ;
        RECT  0.805 1.240 1.065 1.500 ;
        RECT  0.385 1.240 0.805 1.400 ;
        RECT  0.225 0.710 0.385 1.900 ;
        RECT  0.125 0.710 0.225 0.970 ;
        RECT  0.125 1.740 0.225 1.900 ;
    END
END OAI2B11XLMTH

MACRO OAI2B1X1MTH
    CLASS CORE ;
    FOREIGN OAI2B1X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.730 2.770 2.050 ;
        RECT  2.485 0.730 2.560 0.990 ;
        RECT  2.145 1.890 2.560 2.050 ;
        RECT  1.885 1.890 2.145 2.150 ;
        END
        AntennaDiffArea 0.402 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 1.140 2.380 1.710 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.285 1.225 0.755 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 1.145 1.950 1.710 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.800 -0.130 2.870 0.130 ;
        RECT  1.540 -0.130 1.800 0.965 ;
        RECT  0.725 -0.130 1.540 0.130 ;
        RECT  0.125 -0.130 0.725 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 2.740 2.870 3.000 ;
        RECT  2.460 2.230 2.720 3.000 ;
        RECT  1.175 2.740 2.460 3.000 ;
        RECT  0.915 2.100 1.175 3.000 ;
        RECT  0.000 2.740 0.915 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.120 1.260 1.460 1.520 ;
        RECT  0.960 0.865 1.120 1.920 ;
        RECT  0.880 0.865 0.960 1.025 ;
        RECT  0.535 1.760 0.960 1.920 ;
        RECT  0.620 0.765 0.880 1.025 ;
        RECT  0.275 1.760 0.535 2.020 ;
    END
END OAI2B1X1MTH

MACRO OAI2B1X2MTH
    CLASS CORE ;
    FOREIGN OAI2B1X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.355 2.770 2.075 ;
        RECT  2.485 0.355 2.560 0.955 ;
        RECT  2.110 1.915 2.560 2.075 ;
        RECT  1.850 1.915 2.110 2.515 ;
        END
        AntennaDiffArea 0.581 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.130 1.135 2.380 1.735 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.245 1.230 0.720 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 1.135 1.950 1.735 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.725 -0.130 2.870 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 2.740 2.870 3.000 ;
        RECT  2.400 2.315 2.660 3.000 ;
        RECT  1.250 2.740 2.400 3.000 ;
        RECT  0.990 2.145 1.250 3.000 ;
        RECT  0.735 2.740 0.990 3.000 ;
        RECT  0.475 2.570 0.735 3.000 ;
        RECT  0.000 2.740 0.475 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.975 0.355 2.235 0.955 ;
        RECT  1.020 0.355 1.975 0.615 ;
        RECT  1.105 1.230 1.460 1.490 ;
        RECT  0.945 0.815 1.105 1.920 ;
        RECT  0.540 0.815 0.945 0.975 ;
        RECT  0.285 1.760 0.945 1.920 ;
    END
END OAI2B1X2MTH

MACRO OAI2B1X4MTH
    CLASS CORE ;
    FOREIGN OAI2B1X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.955 1.290 4.000 1.940 ;
        RECT  3.775 0.815 3.955 1.940 ;
        RECT  3.615 0.815 3.775 1.045 ;
        RECT  3.765 1.760 3.775 1.940 ;
        RECT  3.505 1.760 3.765 2.400 ;
        RECT  2.340 2.060 3.505 2.240 ;
        RECT  2.080 2.060 2.340 2.320 ;
        END
        AntennaDiffArea 0.974 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.225 3.595 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.260 1.075 1.540 ;
        END
        AntennaGateArea 0.1755 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.925 1.205 2.525 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.845 -0.130 4.510 0.130 ;
        RECT  2.585 -0.130 2.845 0.680 ;
        RECT  0.385 -0.130 2.585 0.130 ;
        RECT  0.125 -0.130 0.385 0.870 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.305 2.740 4.510 3.000 ;
        RECT  4.045 2.115 4.305 3.000 ;
        RECT  3.225 2.740 4.045 3.000 ;
        RECT  2.965 2.420 3.225 3.000 ;
        RECT  1.455 2.740 2.965 3.000 ;
        RECT  1.195 2.230 1.455 3.000 ;
        RECT  0.405 2.740 1.195 3.000 ;
        RECT  0.145 2.570 0.405 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.135 0.385 4.385 0.985 ;
        RECT  3.365 0.385 4.135 0.545 ;
        RECT  3.105 0.385 3.365 1.020 ;
        RECT  2.325 0.860 3.105 1.020 ;
        RECT  2.915 1.200 3.015 1.460 ;
        RECT  2.755 1.200 2.915 1.880 ;
        RECT  1.615 1.720 2.755 1.880 ;
        RECT  2.065 0.385 2.325 1.020 ;
        RECT  1.375 0.580 2.065 0.740 ;
        RECT  1.455 0.920 1.615 1.880 ;
        RECT  0.895 0.920 1.455 1.080 ;
        RECT  0.915 1.720 1.455 1.880 ;
        RECT  1.115 0.355 1.375 0.740 ;
        RECT  0.655 1.720 0.915 2.335 ;
        RECT  0.635 0.765 0.895 1.080 ;
    END
END OAI2B1X4MTH

MACRO OAI2B1X8MTH
    CLASS CORE ;
    FOREIGN OAI2B1X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.150 0.785 7.565 2.395 ;
        RECT  7.070 0.785 7.150 2.140 ;
        RECT  6.285 0.785 7.070 1.115 ;
        RECT  6.505 1.800 7.070 2.140 ;
        RECT  6.165 1.800 6.505 2.440 ;
        RECT  2.765 2.100 6.165 2.440 ;
        END
        AntennaDiffArea 2.084 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.120 1.315 6.720 1.575 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.220 1.100 1.540 ;
        END
        AntennaGateArea 0.351 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.585 1.265 5.135 1.525 ;
        RECT  4.425 0.910 4.585 1.525 ;
        RECT  3.320 0.910 4.425 1.070 ;
        RECT  3.160 0.910 3.320 1.540 ;
        RECT  2.520 1.185 3.160 1.540 ;
        END
        AntennaGateArea 0.8216 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.470 -0.130 8.200 0.130 ;
        RECT  4.210 -0.130 4.470 0.315 ;
        RECT  2.400 -0.130 4.210 0.130 ;
        RECT  2.140 -0.130 2.400 0.645 ;
        RECT  0.385 -0.130 2.140 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.045 2.740 8.200 3.000 ;
        RECT  7.785 1.800 8.045 3.000 ;
        RECT  6.965 2.740 7.785 3.000 ;
        RECT  6.705 2.320 6.965 3.000 ;
        RECT  3.995 2.740 6.705 3.000 ;
        RECT  3.735 2.620 3.995 3.000 ;
        RECT  2.105 2.740 3.735 3.000 ;
        RECT  1.505 2.100 2.105 3.000 ;
        RECT  0.685 2.740 1.505 3.000 ;
        RECT  0.425 1.800 0.685 3.000 ;
        RECT  0.000 2.740 0.425 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.815 0.405 8.075 1.005 ;
        RECT  6.035 0.405 7.815 0.565 ;
        RECT  5.775 0.405 6.035 1.005 ;
        RECT  5.025 0.405 5.775 0.565 ;
        RECT  5.585 1.230 5.775 1.490 ;
        RECT  5.425 1.230 5.585 1.880 ;
        RECT  4.100 1.720 5.425 1.880 ;
        RECT  4.765 0.405 5.025 1.005 ;
        RECT  3.920 0.495 4.765 0.655 ;
        RECT  3.500 1.250 4.100 1.880 ;
        RECT  3.660 0.395 3.920 0.655 ;
        RECT  2.920 0.495 3.660 0.655 ;
        RECT  2.220 1.720 3.500 1.880 ;
        RECT  2.660 0.385 2.920 0.985 ;
        RECT  1.880 0.825 2.660 0.985 ;
        RECT  1.960 1.220 2.220 1.880 ;
        RECT  1.440 1.720 1.960 1.880 ;
        RECT  1.620 0.385 1.880 0.985 ;
        RECT  1.280 0.880 1.440 1.880 ;
        RECT  0.925 0.880 1.280 1.040 ;
        RECT  1.225 1.720 1.280 1.880 ;
        RECT  0.965 1.720 1.225 2.335 ;
        RECT  0.665 0.605 0.925 1.040 ;
    END
END OAI2B1X8MTH

MACRO OAI2B1XLMTH
    CLASS CORE ;
    FOREIGN OAI2B1XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.335 2.770 2.010 ;
        RECT  2.485 0.335 2.560 0.595 ;
        RECT  1.850 1.850 2.560 2.010 ;
        END
        AntennaDiffArea 0.342 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.935 2.380 1.665 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.285 1.225 0.755 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.640 1.205 1.970 1.670 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 -0.130 2.870 0.130 ;
        RECT  1.505 -0.130 1.765 1.025 ;
        RECT  0.725 -0.130 1.505 0.130 ;
        RECT  0.125 -0.130 0.725 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.660 2.740 2.870 3.000 ;
        RECT  2.400 2.195 2.660 3.000 ;
        RECT  2.125 2.740 2.400 3.000 ;
        RECT  1.525 2.570 2.125 3.000 ;
        RECT  1.200 2.740 1.525 3.000 ;
        RECT  0.940 2.105 1.200 3.000 ;
        RECT  0.000 2.740 0.940 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.120 1.260 1.460 1.520 ;
        RECT  0.960 0.865 1.120 1.920 ;
        RECT  0.815 0.865 0.960 1.025 ;
        RECT  0.580 1.760 0.960 1.920 ;
        RECT  0.555 0.765 0.815 1.025 ;
        RECT  0.320 1.760 0.580 2.020 ;
    END
END OAI2B1XLMTH

MACRO OAI2B2X1MTH
    CLASS CORE ;
    FOREIGN OAI2B2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 0.765 2.155 2.100 ;
        RECT  1.565 0.765 1.995 1.130 ;
        RECT  1.465 0.765 1.565 1.025 ;
        END
        AntennaDiffArea 0.582 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.225 3.180 1.640 ;
        RECT  2.690 1.225 2.970 1.560 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.495 1.740 2.810 2.065 ;
        RECT  2.335 1.225 2.495 2.065 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.270 1.225 0.735 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.725 1.310 1.815 1.570 ;
        RECT  1.565 1.310 1.725 1.990 ;
        RECT  1.330 1.700 1.565 1.990 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 3.280 0.130 ;
        RECT  2.485 -0.130 2.745 0.995 ;
        RECT  0.725 -0.130 2.485 0.130 ;
        RECT  0.125 -0.130 0.725 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.215 2.570 3.155 3.000 ;
        RECT  1.825 2.740 2.215 3.000 ;
        RECT  1.145 2.570 1.825 3.000 ;
        RECT  0.885 2.100 1.145 3.000 ;
        RECT  0.000 2.740 0.885 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.105 1.225 1.385 1.485 ;
        RECT  0.945 0.865 1.105 1.920 ;
        RECT  0.815 0.865 0.945 1.025 ;
        RECT  0.285 1.760 0.945 1.920 ;
        RECT  0.555 0.765 0.815 1.025 ;
    END
END OAI2B2X1MTH

MACRO OAI2B2X2MTH
    CLASS CORE ;
    FOREIGN OAI2B2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.800 3.590 2.050 ;
        RECT  1.695 0.800 3.380 0.960 ;
        RECT  2.475 1.890 3.380 2.050 ;
        RECT  2.215 1.890 2.475 2.490 ;
        END
        AntennaDiffArea 0.722 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.950 1.140 3.200 1.710 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 1.140 2.770 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 1.220 0.820 1.575 ;
        END
        AntennaGateArea 0.0871 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.150 2.220 1.665 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.015 -0.130 3.690 0.130 ;
        RECT  2.755 -0.130 3.015 0.270 ;
        RECT  0.735 -0.130 2.755 0.130 ;
        RECT  0.395 -0.130 0.735 0.305 ;
        RECT  0.135 -0.130 0.395 0.985 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.390 2.740 3.690 3.000 ;
        RECT  3.130 2.230 3.390 3.000 ;
        RECT  1.530 2.740 3.130 3.000 ;
        RECT  0.930 2.145 1.530 3.000 ;
        RECT  0.480 2.740 0.930 3.000 ;
        RECT  0.220 2.565 0.480 3.000 ;
        RECT  0.000 2.740 0.220 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.300 0.360 3.560 0.620 ;
        RECT  2.465 0.450 3.300 0.620 ;
        RECT  2.205 0.360 2.465 0.620 ;
        RECT  1.445 0.450 2.205 0.620 ;
        RECT  1.360 1.245 1.555 1.505 ;
        RECT  1.185 0.360 1.445 0.620 ;
        RECT  1.200 0.865 1.360 1.915 ;
        RECT  0.935 0.865 1.200 1.025 ;
        RECT  0.650 1.755 1.200 1.915 ;
        RECT  0.675 0.765 0.935 1.025 ;
        RECT  0.390 1.755 0.650 2.015 ;
    END
END OAI2B2X2MTH

MACRO OAI2B2X4MTH
    CLASS CORE ;
    FOREIGN OAI2B2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.430 0.820 5.640 2.240 ;
        RECT  2.965 0.820 5.430 1.000 ;
        RECT  4.405 2.060 5.430 2.240 ;
        RECT  4.145 2.060 4.405 2.320 ;
        RECT  2.600 2.060 4.145 2.240 ;
        RECT  2.705 0.740 2.965 1.000 ;
        RECT  1.945 0.820 2.705 1.000 ;
        RECT  2.000 2.060 2.600 2.320 ;
        RECT  1.685 0.740 1.945 1.000 ;
        END
        AntennaDiffArea 1.496 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 1.315 5.175 1.575 ;
        RECT  4.915 1.315 5.075 1.880 ;
        RECT  3.755 1.720 4.915 1.880 ;
        RECT  3.380 1.220 3.755 1.880 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 1.220 4.575 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.325 1.245 0.925 1.540 ;
        END
        AntennaGateArea 0.1755 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.195 2.590 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.065 -0.130 5.740 0.130 ;
        RECT  4.805 -0.130 5.065 0.300 ;
        RECT  0.385 -0.130 4.805 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.605 2.740 5.740 3.000 ;
        RECT  5.005 2.420 5.605 3.000 ;
        RECT  3.500 2.740 5.005 3.000 ;
        RECT  3.240 2.420 3.500 3.000 ;
        RECT  1.395 2.740 3.240 3.000 ;
        RECT  0.795 2.100 1.395 3.000 ;
        RECT  0.000 2.740 0.795 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.350 0.380 5.610 0.640 ;
        RECT  4.515 0.480 5.350 0.640 ;
        RECT  4.255 0.380 4.515 0.640 ;
        RECT  3.475 0.480 4.255 0.640 ;
        RECT  3.215 0.380 3.475 0.640 ;
        RECT  2.455 0.380 3.215 0.540 ;
        RECT  3.040 1.220 3.200 1.880 ;
        RECT  1.505 1.720 3.040 1.880 ;
        RECT  2.195 0.380 2.455 0.640 ;
        RECT  1.435 0.380 2.195 0.540 ;
        RECT  1.345 0.905 1.505 1.880 ;
        RECT  1.175 0.380 1.435 0.725 ;
        RECT  0.925 0.905 1.345 1.065 ;
        RECT  0.515 1.720 1.345 1.880 ;
        RECT  0.665 0.620 0.925 1.065 ;
        RECT  0.255 1.720 0.515 2.335 ;
    END
END OAI2B2X4MTH

MACRO OAI2B2X8MTH
    CLASS CORE ;
    FOREIGN OAI2B2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.120 1.495 10.150 2.355 ;
        RECT  9.815 0.770 10.120 2.355 ;
        RECT  6.545 0.770 9.815 0.930 ;
        RECT  2.435 2.060 9.815 2.355 ;
        RECT  6.385 0.745 6.545 0.930 ;
        RECT  2.085 0.745 6.385 0.905 ;
        END
        AntennaDiffArea 2.951 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.585 1.225 9.635 1.485 ;
        RECT  9.425 1.225 9.585 1.880 ;
        RECT  8.275 1.720 9.425 1.880 ;
        RECT  7.675 1.450 8.275 1.880 ;
        RECT  6.235 1.720 7.675 1.880 ;
        RECT  5.840 1.220 6.235 1.880 ;
        END
        AntennaGateArea 0.7982 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.595 1.110 9.195 1.485 ;
        RECT  7.355 1.110 8.595 1.270 ;
        RECT  6.415 1.110 7.355 1.540 ;
        END
        AntennaGateArea 0.7982 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 1.100 1.540 ;
        END
        AntennaGateArea 0.351 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.625 1.225 5.065 1.485 ;
        RECT  4.465 1.085 4.625 1.485 ;
        RECT  3.225 1.085 4.465 1.245 ;
        RECT  2.285 1.085 3.225 1.540 ;
        END
        AntennaGateArea 0.806 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.575 -0.130 10.250 0.130 ;
        RECT  9.315 -0.130 9.575 0.250 ;
        RECT  7.465 -0.130 9.315 0.130 ;
        RECT  7.205 -0.130 7.465 0.250 ;
        RECT  0.385 -0.130 7.205 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.895 2.740 10.250 3.000 ;
        RECT  9.635 2.540 9.895 3.000 ;
        RECT  8.100 2.740 9.635 3.000 ;
        RECT  7.840 2.540 8.100 3.000 ;
        RECT  5.885 2.740 7.840 3.000 ;
        RECT  5.625 2.540 5.885 3.000 ;
        RECT  3.980 2.740 5.625 3.000 ;
        RECT  3.720 2.540 3.980 3.000 ;
        RECT  1.830 2.740 3.720 3.000 ;
        RECT  1.230 2.170 1.830 3.000 ;
        RECT  0.385 2.740 1.230 3.000 ;
        RECT  0.125 1.730 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.915 0.430 10.125 0.590 ;
        RECT  6.655 0.405 6.915 0.590 ;
        RECT  1.785 0.405 6.655 0.565 ;
        RECT  5.315 1.225 5.575 1.880 ;
        RECT  4.135 1.720 5.315 1.880 ;
        RECT  3.535 1.425 4.135 1.880 ;
        RECT  2.065 1.720 3.535 1.880 ;
        RECT  1.805 1.225 2.065 1.880 ;
        RECT  1.445 1.720 1.805 1.880 ;
        RECT  1.625 0.405 1.785 1.025 ;
        RECT  1.285 0.870 1.445 1.880 ;
        RECT  0.925 0.870 1.285 1.030 ;
        RECT  0.925 1.720 1.285 1.880 ;
        RECT  0.665 0.610 0.925 1.030 ;
        RECT  0.665 1.720 0.925 2.330 ;
    END
END OAI2B2X8MTH

MACRO OAI2B2XLMTH
    CLASS CORE ;
    FOREIGN OAI2B2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.995 0.815 2.155 1.975 ;
        RECT  1.500 0.815 1.995 1.130 ;
        END
        AntennaDiffArea 0.376 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 1.225 3.180 1.620 ;
        RECT  2.690 1.225 2.970 1.560 ;
        END
        AntennaGateArea 0.0858 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.495 1.740 2.810 1.950 ;
        RECT  2.335 1.205 2.495 1.950 ;
        END
        AntennaGateArea 0.0858 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.270 1.225 0.735 1.580 ;
        END
        AntennaGateArea 0.0546 ;
    END A1N
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.655 1.310 1.815 1.990 ;
        RECT  1.330 1.700 1.655 1.990 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 -0.130 3.280 0.130 ;
        RECT  2.485 -0.130 2.745 1.025 ;
        RECT  0.725 -0.130 2.485 0.130 ;
        RECT  0.125 -0.130 0.725 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.215 2.570 3.155 3.000 ;
        RECT  1.820 2.740 2.215 3.000 ;
        RECT  1.140 2.570 1.820 3.000 ;
        RECT  0.880 2.230 1.140 3.000 ;
        RECT  0.545 2.740 0.880 3.000 ;
        RECT  0.285 2.610 0.545 3.000 ;
        RECT  0.000 2.740 0.285 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.050 0.310 1.570 0.630 ;
        RECT  1.105 1.240 1.335 1.500 ;
        RECT  0.945 0.815 1.105 1.920 ;
        RECT  0.555 0.815 0.945 0.975 ;
        RECT  0.285 1.760 0.945 1.920 ;
    END
END OAI2B2XLMTH

MACRO OAI2BB1X1MTH
    CLASS CORE ;
    FOREIGN OAI2BB1X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.735 2.360 2.025 ;
        RECT  1.930 0.735 2.150 0.995 ;
        RECT  1.810 1.865 2.150 2.025 ;
        RECT  1.550 1.865 1.810 2.125 ;
        END
        AntennaDiffArea 0.36 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 0.880 1.615 1.345 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.565 0.425 1.130 0.760 ;
        RECT  0.330 0.425 0.565 0.585 ;
        END
        AntennaGateArea 0.0598 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 2.125 1.175 2.360 ;
        END
        AntennaGateArea 0.0598 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 -0.130 2.460 0.130 ;
        RECT  1.260 -0.130 2.200 0.300 ;
        RECT  0.000 -0.130 1.260 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.300 2.740 2.460 3.000 ;
        RECT  1.360 2.565 2.300 3.000 ;
        RECT  1.070 2.740 1.360 3.000 ;
        RECT  0.130 2.565 1.070 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.810 1.225 1.970 1.685 ;
        RECT  0.820 1.525 1.810 1.685 ;
        RECT  0.560 1.525 0.820 1.945 ;
        RECT  0.385 1.525 0.560 1.685 ;
        RECT  0.225 0.765 0.385 1.685 ;
        RECT  0.125 0.765 0.225 1.025 ;
    END
END OAI2BB1X1MTH

MACRO OAI2BB1X2MTH
    CLASS CORE ;
    FOREIGN OAI2BB1X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.310 1.700 2.360 2.125 ;
        RECT  2.150 0.385 2.310 2.125 ;
        RECT  1.930 0.385 2.150 0.985 ;
        RECT  1.880 1.965 2.150 2.125 ;
        RECT  1.620 1.965 1.880 2.465 ;
        END
        AntennaDiffArea 0.571 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 0.880 1.610 1.435 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.855 0.880 1.130 1.170 ;
        RECT  0.650 0.320 0.855 1.170 ;
        RECT  0.330 0.320 0.650 0.555 ;
        END
        AntennaGateArea 0.0975 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 2.110 1.035 2.405 ;
        END
        AntennaGateArea 0.0975 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.305 -0.130 2.460 0.130 ;
        RECT  1.045 -0.130 1.305 0.640 ;
        RECT  0.000 -0.130 1.045 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 2.740 2.460 3.000 ;
        RECT  0.220 2.620 1.160 3.000 ;
        RECT  0.000 2.740 0.220 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.810 1.175 1.970 1.775 ;
        RECT  0.850 1.615 1.810 1.775 ;
        RECT  0.590 1.615 0.850 1.930 ;
        RECT  0.370 1.615 0.590 1.775 ;
        RECT  0.210 0.765 0.370 1.775 ;
    END
END OAI2BB1X2MTH

MACRO OAI2BB1X4MTH
    CLASS CORE ;
    FOREIGN OAI2BB1X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.765 0.405 4.000 2.050 ;
        RECT  2.695 0.405 3.765 0.585 ;
        RECT  3.435 1.870 3.765 2.050 ;
        RECT  3.175 1.870 3.435 2.470 ;
        RECT  2.305 2.060 3.175 2.240 ;
        RECT  2.045 2.060 2.305 2.320 ;
        END
        AntennaDiffArea 1.152 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.695 1.245 2.400 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.165 0.400 1.695 ;
        END
        AntennaGateArea 0.1898 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.165 1.175 1.695 ;
        END
        AntennaGateArea 0.1898 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.445 -0.130 4.100 0.130 ;
        RECT  2.185 -0.130 2.445 0.590 ;
        RECT  1.305 -0.130 2.185 0.130 ;
        RECT  1.045 -0.130 1.305 0.645 ;
        RECT  0.000 -0.130 1.045 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 2.740 4.100 3.000 ;
        RECT  3.715 2.230 3.975 3.000 ;
        RECT  2.875 2.740 3.715 3.000 ;
        RECT  2.615 2.420 2.875 3.000 ;
        RECT  1.735 2.740 2.615 3.000 ;
        RECT  1.235 2.170 1.735 3.000 ;
        RECT  0.385 2.740 1.235 3.000 ;
        RECT  0.125 1.875 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.955 1.225 3.585 1.485 ;
        RECT  1.895 0.770 3.465 0.930 ;
        RECT  2.795 1.225 2.955 1.880 ;
        RECT  1.515 1.720 2.795 1.880 ;
        RECT  1.735 0.430 1.895 0.930 ;
        RECT  1.635 0.430 1.735 0.690 ;
        RECT  1.355 0.825 1.515 1.880 ;
        RECT  0.740 0.825 1.355 0.985 ;
        RECT  0.740 1.875 0.925 2.475 ;
        RECT  0.580 0.825 0.740 2.475 ;
        RECT  0.415 0.825 0.580 0.985 ;
        RECT  0.155 0.385 0.415 0.985 ;
    END
END OAI2BB1X4MTH

MACRO OAI2BB1XLMTH
    CLASS CORE ;
    FOREIGN OAI2BB1XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.765 2.360 2.025 ;
        RECT  1.960 0.765 2.150 1.025 ;
        RECT  1.580 1.865 2.150 2.025 ;
        END
        AntennaDiffArea 0.263 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 0.880 1.615 1.345 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.615 0.375 1.130 0.760 ;
        RECT  0.330 0.375 0.615 0.585 ;
        END
        AntennaGateArea 0.0533 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.355 2.145 1.220 2.360 ;
        END
        AntennaGateArea 0.0533 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 -0.130 2.460 0.130 ;
        RECT  1.295 -0.130 2.235 0.300 ;
        RECT  0.000 -0.130 1.295 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 2.740 2.460 3.000 ;
        RECT  1.395 2.570 2.335 3.000 ;
        RECT  1.070 2.740 1.395 3.000 ;
        RECT  0.130 2.590 1.070 3.000 ;
        RECT  0.000 2.740 0.130 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.810 1.245 1.970 1.685 ;
        RECT  0.820 1.525 1.810 1.685 ;
        RECT  0.560 1.525 0.820 1.965 ;
        RECT  0.385 1.525 0.560 1.685 ;
        RECT  0.225 0.765 0.385 1.685 ;
        RECT  0.125 0.765 0.225 1.025 ;
    END
END OAI2BB1XLMTH

MACRO OAI2BB2X1MTH
    CLASS CORE ;
    FOREIGN OAI2BB2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.610 0.735 2.770 2.400 ;
        RECT  2.485 0.735 2.610 0.995 ;
        RECT  2.105 2.105 2.610 2.400 ;
        END
        AntennaDiffArea 0.42 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.240 1.560 1.810 ;
        END
        AntennaGateArea 0.1235 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.175 2.090 1.585 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.240 1.130 1.735 ;
        RECT  0.830 1.335 0.875 1.735 ;
        END
        AntennaGateArea 0.0598 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 0.675 0.355 0.935 ;
        RECT  0.100 0.675 0.310 1.335 ;
        END
        AntennaGateArea 0.0598 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 -0.130 2.870 0.130 ;
        RECT  1.565 -0.130 1.825 0.415 ;
        RECT  0.355 -0.130 1.565 0.130 ;
        RECT  0.125 -0.130 0.355 0.495 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 2.740 2.870 3.000 ;
        RECT  2.485 2.580 2.745 3.000 ;
        RECT  1.355 2.740 2.485 3.000 ;
        RECT  0.855 2.425 1.355 3.000 ;
        RECT  0.675 2.740 0.855 3.000 ;
        RECT  0.175 2.425 0.675 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.270 1.290 2.430 1.925 ;
        RECT  1.925 1.765 2.270 1.925 ;
        RECT  1.975 0.735 2.235 0.995 ;
        RECT  1.280 0.835 1.975 0.995 ;
        RECT  1.765 1.765 1.925 2.170 ;
        RECT  0.840 2.010 1.765 2.170 ;
        RECT  1.020 0.835 1.280 1.060 ;
        RECT  0.695 0.355 1.275 0.515 ;
        RECT  0.650 1.915 0.840 2.170 ;
        RECT  0.650 0.355 0.695 1.215 ;
        RECT  0.535 0.355 0.650 2.170 ;
        RECT  0.490 1.055 0.535 2.170 ;
    END
END OAI2BB2X1MTH

MACRO OAI2BB2X2MTH
    CLASS CORE ;
    FOREIGN OAI2BB2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.945 0.410 3.180 1.925 ;
        RECT  2.560 1.765 2.945 1.925 ;
        RECT  2.300 1.765 2.560 2.395 ;
        END
        AntennaDiffArea 0.667 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.180 1.805 1.585 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 1.175 2.420 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.175 1.150 1.625 ;
        END
        AntennaGateArea 0.0962 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.980 0.355 1.580 ;
        END
        AntennaGateArea 0.0962 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.065 -0.130 3.280 0.130 ;
        RECT  0.125 -0.130 1.065 0.405 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 2.740 3.280 3.000 ;
        RECT  2.895 2.105 3.155 3.000 ;
        RECT  1.565 2.740 2.895 3.000 ;
        RECT  1.305 1.765 1.565 3.000 ;
        RECT  0.940 2.740 1.305 3.000 ;
        RECT  0.680 2.540 0.940 3.000 ;
        RECT  0.335 2.740 0.680 3.000 ;
        RECT  0.135 1.760 0.335 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.605 0.835 2.765 1.485 ;
        RECT  1.395 0.395 2.645 0.655 ;
        RECT  1.145 0.835 2.605 0.995 ;
        RECT  0.885 0.735 1.145 0.995 ;
        RECT  0.695 1.805 0.940 2.000 ;
        RECT  0.695 0.835 0.885 0.995 ;
        RECT  0.535 0.835 0.695 2.000 ;
    END
END OAI2BB2X2MTH

MACRO OAI2BB2X4MTH
    CLASS CORE ;
    FOREIGN OAI2BB2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 1.765 3.705 2.405 ;
        RECT  2.360 1.765 3.445 1.925 ;
        RECT  2.235 1.290 2.360 1.925 ;
        RECT  2.075 0.735 2.235 1.925 ;
        RECT  1.975 0.735 2.075 0.995 ;
        RECT  1.990 1.765 2.075 1.925 ;
        RECT  1.730 1.765 1.990 2.405 ;
        END
        AntennaDiffArea 0.952 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.305 1.245 4.405 1.505 ;
        RECT  4.145 0.985 4.305 1.505 ;
        RECT  3.085 0.985 4.145 1.145 ;
        RECT  2.925 0.985 3.085 1.585 ;
        RECT  2.560 1.235 2.925 1.585 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.275 1.325 3.875 1.585 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.245 1.350 1.585 ;
        END
        AntennaGateArea 0.1885 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.085 0.385 1.655 ;
        END
        AntennaGateArea 0.1885 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.245 -0.130 4.920 0.130 ;
        RECT  3.985 -0.130 4.245 0.460 ;
        RECT  0.385 -0.130 3.985 0.130 ;
        RECT  0.125 -0.130 0.385 0.905 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.565 2.740 4.920 3.000 ;
        RECT  4.305 1.765 4.565 3.000 ;
        RECT  2.845 2.740 4.305 3.000 ;
        RECT  2.245 2.115 2.845 3.000 ;
        RECT  1.445 2.740 2.245 3.000 ;
        RECT  1.185 1.765 1.445 3.000 ;
        RECT  0.385 2.740 1.185 3.000 ;
        RECT  0.125 1.835 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.535 0.385 4.795 0.985 ;
        RECT  3.695 0.640 4.535 0.800 ;
        RECT  3.435 0.540 3.695 0.800 ;
        RECT  2.745 0.640 3.435 0.800 ;
        RECT  2.485 0.395 2.745 0.995 ;
        RECT  1.725 0.395 2.485 0.555 ;
        RECT  1.715 1.235 1.815 1.495 ;
        RECT  1.465 0.395 1.725 0.720 ;
        RECT  1.555 0.900 1.715 1.495 ;
        RECT  1.215 0.900 1.555 1.060 ;
        RECT  0.955 0.385 1.215 1.060 ;
        RECT  0.725 0.900 0.955 1.060 ;
        RECT  0.725 1.765 0.905 2.365 ;
        RECT  0.565 0.900 0.725 2.365 ;
    END
END OAI2BB2X4MTH

MACRO OAI2BB2X8MTH
    CLASS CORE ;
    FOREIGN OAI2BB2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.205 1.905 7.465 2.505 ;
        RECT  5.600 1.905 7.205 2.255 ;
        RECT  5.340 1.905 5.600 2.505 ;
        RECT  5.160 1.905 5.340 2.255 ;
        RECT  4.810 1.665 5.160 2.255 ;
        RECT  4.105 1.665 4.810 2.015 ;
        RECT  4.045 0.745 4.105 2.015 ;
        RECT  3.785 0.745 4.045 2.405 ;
        RECT  3.705 0.745 3.785 2.015 ;
        RECT  2.825 0.745 3.705 1.065 ;
        RECT  2.965 1.665 3.705 2.015 ;
        RECT  2.705 1.665 2.965 2.405 ;
        END
        AntennaDiffArea 1.956 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.065 1.245 8.205 1.505 ;
        RECT  7.905 0.985 8.065 1.505 ;
        RECT  6.725 0.985 7.905 1.145 ;
        RECT  6.120 0.985 6.725 1.345 ;
        RECT  6.075 0.985 6.120 1.145 ;
        RECT  5.915 0.920 6.075 1.145 ;
        RECT  4.895 0.920 5.915 1.080 ;
        RECT  4.570 0.920 4.895 1.445 ;
        END
        AntennaGateArea 0.8216 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.035 1.330 7.635 1.685 ;
        RECT  5.825 1.525 7.035 1.685 ;
        RECT  5.390 1.305 5.825 1.685 ;
        RECT  5.225 1.305 5.390 1.495 ;
        END
        AntennaGateArea 0.8216 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 1.245 2.005 1.580 ;
        RECT  1.555 0.885 1.715 1.580 ;
        RECT  0.695 0.885 1.555 1.045 ;
        RECT  0.535 0.885 0.695 1.505 ;
        RECT  0.295 1.245 0.535 1.505 ;
        END
        AntennaGateArea 0.377 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.225 1.375 1.580 ;
        END
        AntennaGateArea 0.377 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.015 -0.130 8.610 0.130 ;
        RECT  6.755 -0.130 7.015 0.460 ;
        RECT  1.245 -0.130 6.755 0.130 ;
        RECT  0.985 -0.130 1.245 0.365 ;
        RECT  0.000 -0.130 0.985 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.325 2.740 8.610 3.000 ;
        RECT  8.065 1.795 8.325 3.000 ;
        RECT  6.560 2.740 8.065 3.000 ;
        RECT  6.300 2.435 6.560 3.000 ;
        RECT  4.630 2.740 6.300 3.000 ;
        RECT  4.370 2.195 4.630 3.000 ;
        RECT  3.505 2.740 4.370 3.000 ;
        RECT  3.245 2.195 3.505 3.000 ;
        RECT  2.425 2.740 3.245 3.000 ;
        RECT  2.165 2.105 2.425 3.000 ;
        RECT  0.385 2.740 2.165 3.000 ;
        RECT  0.125 1.755 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.245 0.365 8.490 0.965 ;
        RECT  7.555 0.645 8.245 0.805 ;
        RECT  7.295 0.480 7.555 0.805 ;
        RECT  6.475 0.645 7.295 0.805 ;
        RECT  6.215 0.355 6.475 0.805 ;
        RECT  5.545 0.355 6.215 0.515 ;
        RECT  5.285 0.355 5.545 0.740 ;
        RECT  4.615 0.355 5.285 0.515 ;
        RECT  4.355 0.355 4.615 0.690 ;
        RECT  3.595 0.355 4.355 0.515 ;
        RECT  3.335 0.355 3.595 0.565 ;
        RECT  2.425 1.285 3.525 1.445 ;
        RECT  2.285 0.355 3.335 0.515 ;
        RECT  2.265 0.900 2.425 1.925 ;
        RECT  2.055 0.900 2.265 1.060 ;
        RECT  1.885 1.765 2.265 1.925 ;
        RECT  1.895 0.545 2.055 1.060 ;
        RECT  0.355 0.545 1.895 0.705 ;
        RECT  1.625 1.765 1.885 2.365 ;
        RECT  0.925 1.765 1.625 1.925 ;
        RECT  0.665 1.765 0.925 2.365 ;
        RECT  0.125 0.380 0.355 0.980 ;
    END
END OAI2BB2X8MTH

MACRO OAI2BB2XLMTH
    CLASS CORE ;
    FOREIGN OAI2BB2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.755 2.770 1.955 ;
        RECT  2.485 0.755 2.560 1.015 ;
        RECT  2.295 1.795 2.560 1.955 ;
        RECT  2.135 1.795 2.295 2.055 ;
        END
        AntennaDiffArea 0.268 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.455 1.090 1.615 1.590 ;
        RECT  1.330 1.230 1.455 1.590 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 2.275 2.095 2.560 ;
        RECT  1.670 2.110 1.960 2.560 ;
        END
        AntennaGateArea 0.0858 ;
    END B0
    PIN A1N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.235 1.150 1.685 ;
        END
        AntennaGateArea 0.0533 ;
    END A1N
    PIN A0N
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.355 1.695 ;
        END
        AntennaGateArea 0.0533 ;
    END A0N
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.495 -0.130 2.870 0.130 ;
        RECT  1.555 -0.130 2.495 0.405 ;
        RECT  0.000 -0.130 1.555 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 2.740 2.870 3.000 ;
        RECT  2.485 2.405 2.745 3.000 ;
        RECT  1.355 2.740 2.485 3.000 ;
        RECT  0.855 2.365 1.355 3.000 ;
        RECT  0.675 2.740 0.855 3.000 ;
        RECT  0.175 2.365 0.675 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.220 1.355 2.380 1.615 ;
        RECT  1.975 0.750 2.235 1.015 ;
        RECT  1.955 1.455 2.220 1.615 ;
        RECT  1.235 0.750 1.975 0.910 ;
        RECT  1.795 1.455 1.955 1.930 ;
        RECT  1.490 1.770 1.795 1.930 ;
        RECT  1.330 1.770 1.490 2.055 ;
        RECT  0.695 1.895 1.330 2.055 ;
        RECT  0.695 0.355 1.235 0.515 ;
        RECT  0.975 0.750 1.235 1.055 ;
        RECT  0.535 0.355 0.695 2.055 ;
    END
END OAI2BB2XLMTH

MACRO OAI31X1MTH
    CLASS CORE ;
    FOREIGN OAI31X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.675 2.360 1.990 ;
        RECT  2.075 0.675 2.200 0.935 ;
        RECT  2.150 1.700 2.200 1.990 ;
        RECT  1.695 1.830 2.150 1.990 ;
        RECT  1.435 1.830 1.695 2.090 ;
        END
        AntennaDiffArea 0.358 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.095 1.985 1.625 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.180 0.455 1.560 ;
        RECT  0.100 1.180 0.310 1.620 ;
        END
        AntennaGateArea 0.1274 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.075 0.995 1.950 ;
        RECT  0.470 1.740 0.835 1.950 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.265 1.095 1.545 1.650 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 -0.130 2.460 0.130 ;
        RECT  0.220 -0.130 1.160 0.345 ;
        RECT  0.000 -0.130 0.220 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.235 2.740 2.460 3.000 ;
        RECT  1.975 2.170 2.235 3.000 ;
        RECT  0.385 2.740 1.975 3.000 ;
        RECT  0.125 2.110 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.570 0.725 1.825 0.885 ;
    END
END OAI31X1MTH

MACRO OAI31X2MTH
    CLASS CORE ;
    FOREIGN OAI31X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.380 2.770 1.990 ;
        RECT  2.395 0.380 2.560 0.980 ;
        RECT  1.930 1.780 2.560 1.990 ;
        RECT  1.670 1.780 1.930 2.405 ;
        END
        AntennaDiffArea 0.571 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.055 1.165 2.380 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.350 1.225 0.740 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.300 1.230 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.120 1.760 1.485 ;
        RECT  1.480 0.920 1.700 1.485 ;
        RECT  1.290 0.920 1.480 1.130 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.580 -0.130 2.870 0.130 ;
        RECT  1.320 -0.130 1.580 0.400 ;
        RECT  0.480 -0.130 1.320 0.130 ;
        RECT  0.220 -0.130 0.480 1.025 ;
        RECT  0.000 -0.130 0.220 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.470 2.740 2.870 3.000 ;
        RECT  2.210 2.170 2.470 3.000 ;
        RECT  0.590 2.740 2.210 3.000 ;
        RECT  0.330 1.760 0.590 3.000 ;
        RECT  0.000 2.740 0.330 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.880 0.385 2.140 0.985 ;
        RECT  1.030 0.580 1.880 0.740 ;
        RECT  0.770 0.385 1.030 0.985 ;
    END
END OAI31X2MTH

MACRO OAI31X4MTH
    CLASS CORE ;
    FOREIGN OAI31X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 0.835 4.420 1.990 ;
        RECT  3.875 0.835 4.200 1.015 ;
        RECT  3.805 1.810 4.200 1.990 ;
        RECT  3.615 0.735 3.875 1.015 ;
        RECT  3.625 1.810 3.805 2.485 ;
        RECT  1.685 2.305 3.625 2.485 ;
        END
        AntennaDiffArea 0.912 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 1.225 4.015 1.485 ;
        RECT  3.380 1.225 3.590 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.975 1.410 3.075 1.570 ;
        RECT  2.815 1.410 2.975 2.125 ;
        RECT  0.720 1.965 2.815 2.125 ;
        RECT  0.560 1.290 0.720 2.125 ;
        RECT  0.445 1.290 0.560 1.580 ;
        END
        AntennaGateArea 0.3978 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.495 1.415 2.595 1.575 ;
        RECT  2.335 1.415 2.495 1.785 ;
        RECT  1.215 1.625 2.335 1.785 ;
        RECT  0.920 1.290 1.215 1.785 ;
        END
        AntennaGateArea 0.3978 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.990 1.130 2.115 1.445 ;
        RECT  1.700 0.920 1.990 1.445 ;
        RECT  1.515 1.130 1.700 1.445 ;
        END
        AntennaGateArea 0.3978 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 -0.130 4.510 0.130 ;
        RECT  2.565 -0.130 2.825 0.565 ;
        RECT  0.000 -0.130 2.565 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 2.420 4.385 3.000 ;
        RECT  0.380 2.740 4.125 3.000 ;
        RECT  0.135 1.760 0.380 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.125 0.395 4.385 0.655 ;
        RECT  3.365 0.395 4.125 0.555 ;
        RECT  3.265 0.395 3.365 0.775 ;
        RECT  3.105 0.395 3.265 0.905 ;
        RECT  2.330 0.745 3.105 0.905 ;
        RECT  2.170 0.460 2.330 0.905 ;
        RECT  2.025 0.460 2.170 0.740 ;
        RECT  1.335 0.580 2.025 0.740 ;
        RECT  1.075 0.395 1.335 0.995 ;
        RECT  0.390 0.580 1.075 0.740 ;
        RECT  0.130 0.395 0.390 0.995 ;
    END
END OAI31X4MTH

MACRO OAI31XLMTH
    CLASS CORE ;
    FOREIGN OAI31XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.200 0.355 2.360 1.990 ;
        RECT  2.075 0.355 2.200 0.515 ;
        RECT  2.150 1.700 2.200 1.990 ;
        RECT  1.475 1.760 2.150 1.990 ;
        END
        AntennaDiffArea 0.359 ;
    END Y
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.725 1.105 1.985 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.180 0.460 1.560 ;
        RECT  0.100 1.180 0.310 1.625 ;
        END
        AntennaGateArea 0.0702 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.945 1.115 1.045 1.375 ;
        RECT  0.785 1.115 0.945 1.950 ;
        RECT  0.470 1.740 0.785 1.950 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.225 1.100 1.545 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.825 -0.130 2.460 0.130 ;
        RECT  1.245 -0.130 1.825 0.345 ;
        RECT  1.065 -0.130 1.245 0.130 ;
        RECT  0.125 -0.130 1.065 0.345 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 2.740 2.460 3.000 ;
        RECT  2.065 2.170 2.325 3.000 ;
        RECT  1.695 2.740 2.065 3.000 ;
        RECT  0.755 2.570 1.695 3.000 ;
        RECT  0.385 2.740 0.755 3.000 ;
        RECT  0.125 2.110 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.595 0.675 1.855 0.925 ;
        RECT  0.830 0.675 1.595 0.835 ;
        RECT  0.570 0.675 0.830 0.935 ;
    END
END OAI31XLMTH

MACRO OAI32X1MTH
    CLASS CORE ;
    FOREIGN OAI32X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.825 2.380 2.400 ;
        RECT  2.175 0.775 2.335 2.400 ;
        RECT  1.975 0.775 2.175 0.935 ;
        RECT  2.150 1.825 2.175 2.400 ;
        RECT  1.545 1.825 2.150 2.085 ;
        END
        AntennaDiffArea 0.49 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.570 1.210 2.770 1.940 ;
        RECT  2.515 1.210 2.570 1.650 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.170 1.995 1.645 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.210 0.565 1.470 ;
        RECT  0.100 0.880 0.310 1.470 ;
        END
        AntennaGateArea 0.1274 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.310 0.995 1.990 ;
        RECT  0.510 1.700 0.835 1.990 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.335 1.210 1.520 1.470 ;
        RECT  1.175 0.920 1.335 1.470 ;
        RECT  0.880 0.920 1.175 1.130 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.325 -0.130 2.870 0.130 ;
        RECT  1.065 -0.130 1.325 0.370 ;
        RECT  0.000 -0.130 1.065 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 2.740 2.870 3.000 ;
        RECT  1.805 2.580 2.745 3.000 ;
        RECT  1.065 2.740 1.805 3.000 ;
        RECT  0.125 2.555 1.065 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.535 0.435 2.695 0.990 ;
        RECT  1.675 0.435 2.535 0.595 ;
        RECT  1.515 0.435 1.675 0.990 ;
        RECT  0.735 0.550 1.515 0.710 ;
        RECT  0.575 0.550 0.735 0.810 ;
    END
END OAI32X1MTH

MACRO OAI32X2MTH
    CLASS CORE ;
    FOREIGN OAI32X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.700 1.700 2.770 1.990 ;
        RECT  2.540 0.710 2.700 1.990 ;
        RECT  2.355 0.710 2.540 0.970 ;
        RECT  1.950 1.810 2.540 1.990 ;
        RECT  1.690 1.810 1.950 2.410 ;
        END
        AntennaDiffArea 0.784 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.960 1.230 3.180 1.845 ;
        RECT  2.880 1.230 2.960 1.490 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.890 1.230 2.360 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.380 1.230 0.655 1.490 ;
        RECT  0.100 0.880 0.380 1.490 ;
        END
        AntennaGateArea 0.2054 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.995 1.310 1.165 1.470 ;
        RECT  0.835 1.310 0.995 1.990 ;
        RECT  0.510 1.700 0.835 1.990 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.440 0.920 1.650 1.490 ;
        RECT  0.880 0.920 1.440 1.130 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 -0.130 3.280 0.130 ;
        RECT  1.305 -0.130 1.565 0.400 ;
        RECT  0.475 -0.130 1.305 0.130 ;
        RECT  0.215 -0.130 0.475 0.700 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.970 2.740 3.280 3.000 ;
        RECT  2.710 2.170 2.970 3.000 ;
        RECT  0.475 2.740 2.710 3.000 ;
        RECT  0.215 2.170 0.475 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.880 0.365 3.140 0.980 ;
        RECT  2.105 0.365 2.880 0.525 ;
        RECT  1.845 0.365 2.105 0.980 ;
        RECT  1.025 0.580 1.845 0.740 ;
        RECT  0.765 0.480 1.025 0.740 ;
    END
END OAI32X2MTH

MACRO OAI32X4MTH
    CLASS CORE ;
    FOREIGN OAI32X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.430 0.785 5.640 2.360 ;
        RECT  3.825 0.785 5.430 0.965 ;
        RECT  4.595 2.180 5.430 2.360 ;
        RECT  4.335 2.100 4.595 2.360 ;
        RECT  1.925 2.180 4.335 2.360 ;
        RECT  1.665 2.100 1.925 2.360 ;
        END
        AntennaDiffArea 1.27 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.150 1.230 5.250 1.490 ;
        RECT  4.990 1.230 5.150 1.900 ;
        RECT  3.940 1.740 4.990 1.900 ;
        RECT  3.680 1.210 3.940 1.900 ;
        RECT  3.180 1.700 3.680 1.900 ;
        RECT  2.970 1.700 3.180 1.990 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.230 4.765 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.035 1.230 3.180 1.490 ;
        RECT  2.875 0.825 3.035 1.490 ;
        RECT  0.700 0.825 2.875 0.985 ;
        RECT  0.540 0.825 0.700 1.580 ;
        RECT  0.100 1.230 0.540 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.395 1.230 2.655 1.880 ;
        RECT  1.170 1.720 2.395 1.880 ;
        RECT  0.880 1.230 1.170 1.950 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.495 1.260 2.095 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.025 -0.130 5.740 0.130 ;
        RECT  2.765 -0.130 3.025 0.305 ;
        RECT  1.925 -0.130 2.765 0.130 ;
        RECT  1.665 -0.130 1.925 0.305 ;
        RECT  0.000 -0.130 1.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.460 2.740 5.740 3.000 ;
        RECT  5.200 2.540 5.460 3.000 ;
        RECT  3.710 2.740 5.200 3.000 ;
        RECT  3.110 2.540 3.710 3.000 ;
        RECT  0.505 2.740 3.110 3.000 ;
        RECT  0.245 1.790 0.505 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.355 0.405 5.615 0.605 ;
        RECT  4.595 0.445 5.355 0.605 ;
        RECT  4.335 0.405 4.595 0.605 ;
        RECT  3.575 0.445 4.335 0.605 ;
        RECT  3.315 0.445 3.575 0.995 ;
        RECT  2.475 0.485 3.315 0.645 ;
        RECT  2.215 0.385 2.475 0.645 ;
        RECT  1.375 0.485 2.215 0.645 ;
        RECT  1.115 0.385 1.375 0.645 ;
        RECT  0.360 0.485 1.115 0.645 ;
        RECT  0.125 0.380 0.360 0.980 ;
    END
END OAI32X4MTH

MACRO OAI32XLMTH
    CLASS CORE ;
    FOREIGN OAI32XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 1.825 2.360 2.400 ;
        RECT  2.175 0.760 2.335 2.400 ;
        RECT  2.055 0.760 2.175 1.020 ;
        RECT  2.150 1.825 2.175 2.400 ;
        RECT  1.545 1.825 2.150 2.085 ;
        END
        AntennaDiffArea 0.31 ;
    END Y
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 1.210 2.770 1.845 ;
        RECT  2.515 1.210 2.550 1.730 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.190 1.995 1.645 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 0.565 1.465 ;
        RECT  0.100 0.880 0.310 1.465 ;
        END
        AntennaGateArea 0.0702 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.835 1.205 0.995 1.860 ;
        RECT  0.720 1.700 0.835 1.860 ;
        RECT  0.510 1.700 0.720 1.990 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.365 1.255 1.515 1.515 ;
        RECT  1.175 1.255 1.365 2.360 ;
        RECT  0.880 2.150 1.175 2.360 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.315 -0.130 2.870 0.130 ;
        RECT  1.055 -0.130 1.315 1.020 ;
        RECT  0.385 -0.130 1.055 0.130 ;
        RECT  0.125 -0.130 0.385 0.310 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.745 2.740 2.870 3.000 ;
        RECT  1.805 2.580 2.745 3.000 ;
        RECT  1.065 2.740 1.805 3.000 ;
        RECT  0.125 2.540 1.065 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
END OAI32XLMTH

MACRO OAI33X1MTH
    CLASS CORE ;
    FOREIGN OAI33X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.710 3.590 1.920 ;
        RECT  2.225 0.710 3.380 0.870 ;
        RECT  2.745 1.760 3.380 1.920 ;
        RECT  2.585 1.760 2.745 2.290 ;
        RECT  1.760 2.130 2.585 2.290 ;
        RECT  1.500 1.810 1.760 2.290 ;
        END
        AntennaDiffArea 0.53 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.215 0.515 1.560 ;
        RECT  0.100 1.215 0.310 1.640 ;
        END
        AntennaGateArea 0.1274 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.875 1.215 1.035 1.950 ;
        RECT  0.470 1.740 0.875 1.950 ;
        END
        AntennaGateArea 0.1274 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 1.125 1.540 1.595 ;
        END
        AntennaGateArea 0.1274 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.060 3.180 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 1.060 2.625 1.320 ;
        RECT  2.245 1.060 2.405 1.950 ;
        RECT  2.110 1.740 2.245 1.950 ;
        END
        AntennaGateArea 0.1274 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 1.060 2.065 1.320 ;
        RECT  1.740 1.060 2.015 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.425 -0.130 3.690 0.130 ;
        RECT  0.825 -0.130 1.425 0.330 ;
        RECT  0.385 -0.130 0.825 0.130 ;
        RECT  0.125 -0.130 0.385 0.920 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 2.740 3.690 3.000 ;
        RECT  2.925 2.100 3.525 3.000 ;
        RECT  1.090 2.740 2.925 3.000 ;
        RECT  0.150 2.570 1.090 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.975 0.355 3.025 0.515 ;
        RECT  1.815 0.355 1.975 0.875 ;
        RECT  0.645 0.715 1.815 0.875 ;
    END
END OAI33X1MTH

MACRO OAI33X2MTH
    CLASS CORE ;
    FOREIGN OAI33X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.380 3.590 2.085 ;
        RECT  3.305 0.380 3.380 1.020 ;
        RECT  2.905 1.885 3.380 2.085 ;
        RECT  2.485 0.820 3.305 1.020 ;
        RECT  2.705 1.885 2.905 2.410 ;
        RECT  1.855 2.210 2.705 2.410 ;
        RECT  2.225 0.760 2.485 1.020 ;
        RECT  1.595 1.810 1.855 2.410 ;
        END
        AntennaDiffArea 1.051 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.150 0.565 1.505 ;
        RECT  0.100 1.150 0.310 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.825 1.310 1.085 1.950 ;
        RECT  0.470 1.740 0.825 1.950 ;
        END
        AntennaGateArea 0.2054 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.355 0.920 1.515 1.485 ;
        RECT  0.880 0.920 1.355 1.130 ;
        END
        AntennaGateArea 0.2054 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.835 1.205 3.180 1.705 ;
        END
        AntennaGateArea 0.2054 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.525 1.225 2.655 1.485 ;
        RECT  2.275 1.225 2.525 1.950 ;
        RECT  2.110 1.740 2.275 1.950 ;
        END
        AntennaGateArea 0.2054 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.700 1.205 2.095 1.540 ;
        END
        AntennaGateArea 0.2054 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.385 -0.130 3.690 0.130 ;
        RECT  0.125 -0.130 0.385 0.970 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 2.740 3.690 3.000 ;
        RECT  3.085 2.265 3.345 3.000 ;
        RECT  0.385 2.740 3.085 3.000 ;
        RECT  0.125 2.110 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.765 0.320 3.025 0.640 ;
        RECT  1.975 0.320 2.765 0.580 ;
        RECT  1.715 0.320 1.975 0.740 ;
        RECT  0.645 0.480 1.715 0.740 ;
    END
END OAI33X2MTH

MACRO OAI33X4MTH
    CLASS CORE ;
    FOREIGN OAI33X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 0.745 6.870 2.440 ;
        RECT  3.595 0.745 6.660 0.905 ;
        RECT  1.745 2.260 6.660 2.440 ;
        RECT  1.485 2.060 1.745 2.440 ;
        END
        AntennaDiffArea 1.889 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.965 1.230 3.065 1.490 ;
        RECT  2.805 0.770 2.965 1.490 ;
        RECT  0.565 0.770 2.805 0.930 ;
        RECT  0.405 0.770 0.565 1.490 ;
        RECT  0.310 1.150 0.405 1.490 ;
        RECT  0.100 1.150 0.310 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.485 1.230 2.585 1.490 ;
        RECT  2.325 1.230 2.485 1.880 ;
        RECT  1.075 1.720 2.325 1.880 ;
        RECT  0.815 1.230 1.075 1.950 ;
        RECT  0.470 1.740 0.815 1.950 ;
        END
        AntennaGateArea 0.4108 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.260 2.045 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.230 1.230 6.390 2.080 ;
        RECT  3.495 1.920 6.230 2.080 ;
        RECT  3.335 1.230 3.495 2.080 ;
        RECT  2.970 1.700 3.335 2.080 ;
        END
        AntennaGateArea 0.4108 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 1.085 5.640 1.400 ;
        RECT  4.040 1.085 5.380 1.245 ;
        RECT  3.750 1.085 4.040 1.540 ;
        END
        AntennaGateArea 0.4108 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.840 1.290 6.050 1.740 ;
        RECT  5.125 1.580 5.840 1.740 ;
        RECT  4.845 1.425 5.125 1.740 ;
        END
        AntennaGateArea 0.403 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 -0.130 6.970 0.130 ;
        RECT  1.615 -0.130 1.875 0.250 ;
        RECT  0.000 -0.130 1.615 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.705 2.740 6.970 3.000 ;
        RECT  6.105 2.620 6.705 3.000 ;
        RECT  3.275 2.740 6.105 3.000 ;
        RECT  3.015 2.620 3.275 3.000 ;
        RECT  0.385 2.740 3.015 3.000 ;
        RECT  0.125 2.110 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.345 0.405 6.845 0.565 ;
        RECT  3.085 0.405 3.345 0.590 ;
        RECT  0.125 0.430 3.085 0.590 ;
    END
END OAI33X4MTH

MACRO OAI33XLMTH
    CLASS CORE ;
    FOREIGN OAI33XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.380 0.710 3.590 1.920 ;
        RECT  2.165 0.710 3.380 0.870 ;
        RECT  2.745 1.760 3.380 1.920 ;
        RECT  2.585 1.760 2.745 2.290 ;
        RECT  1.760 2.130 2.585 2.290 ;
        RECT  1.500 1.775 1.760 2.290 ;
        END
        AntennaDiffArea 0.378 ;
    END Y
    PIN B2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.215 0.515 1.560 ;
        RECT  0.100 1.215 0.310 1.650 ;
        END
        AntennaGateArea 0.0702 ;
    END B2
    PIN B1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 1.215 1.060 1.950 ;
        RECT  0.470 1.740 0.900 1.950 ;
        END
        AntennaGateArea 0.0702 ;
    END B1
    PIN B0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 1.125 1.540 1.595 ;
        END
        AntennaGateArea 0.0702 ;
    END B0
    PIN A2
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.925 1.060 3.180 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A2
    PIN A1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 1.060 2.625 1.320 ;
        RECT  2.245 1.060 2.405 1.950 ;
        RECT  2.110 1.740 2.245 1.950 ;
        END
        AntennaGateArea 0.0702 ;
    END A1
    PIN A0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.015 1.080 2.065 1.340 ;
        RECT  1.740 1.080 2.015 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END A0
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.505 -0.130 3.690 0.130 ;
        RECT  3.245 -0.130 3.505 0.300 ;
        RECT  1.505 -0.130 3.245 0.130 ;
        RECT  0.905 -0.130 1.505 0.330 ;
        RECT  0.725 -0.130 0.905 0.130 ;
        RECT  0.125 -0.130 0.725 0.330 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.525 2.740 3.690 3.000 ;
        RECT  2.925 2.100 3.525 3.000 ;
        RECT  2.430 2.740 2.925 3.000 ;
        RECT  1.490 2.470 2.430 3.000 ;
        RECT  1.090 2.740 1.490 3.000 ;
        RECT  0.150 2.470 1.090 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.975 0.355 2.995 0.515 ;
        RECT  1.815 0.355 1.975 0.875 ;
        RECT  0.570 0.715 1.815 0.875 ;
    END
END OAI33XLMTH

MACRO OR2X12MTH
    CLASS CORE ;
    FOREIGN OR2X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.635 0.425 6.255 2.440 ;
        RECT  5.065 0.425 5.635 1.135 ;
        RECT  5.045 1.735 5.635 2.440 ;
        RECT  4.255 0.745 5.065 1.135 ;
        RECT  4.285 1.735 5.045 2.125 ;
        RECT  4.025 1.735 4.285 2.440 ;
        RECT  4.095 0.425 4.255 1.135 ;
        END
        AntennaDiffArea 1.832 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.480 1.225 3.575 1.485 ;
        RECT  3.320 1.225 3.480 2.440 ;
        RECT  2.360 2.280 3.320 2.440 ;
        RECT  1.910 2.110 2.360 2.440 ;
        RECT  1.740 1.225 1.910 2.440 ;
        RECT  0.685 2.280 1.740 2.440 ;
        RECT  0.525 1.225 0.685 2.440 ;
        RECT  0.385 1.225 0.525 1.485 ;
        END
        AntennaGateArea 0.637 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.590 1.225 2.750 1.485 ;
        RECT  2.255 1.225 2.590 1.385 ;
        RECT  2.095 0.880 2.255 1.385 ;
        RECT  1.540 0.880 2.095 1.040 ;
        RECT  1.205 0.880 1.540 1.545 ;
        END
        AntennaGateArea 0.637 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.840 -0.130 6.970 0.130 ;
        RECT  6.580 -0.130 6.840 0.980 ;
        RECT  4.815 -0.130 6.580 0.130 ;
        RECT  4.555 -0.130 4.815 0.565 ;
        RECT  3.725 -0.130 4.555 0.130 ;
        RECT  3.465 -0.130 3.725 0.655 ;
        RECT  3.205 -0.130 3.465 0.130 ;
        RECT  2.945 -0.130 3.205 0.640 ;
        RECT  2.105 -0.130 2.945 0.130 ;
        RECT  1.845 -0.130 2.105 0.360 ;
        RECT  0.685 -0.130 1.845 0.130 ;
        RECT  0.445 -0.130 0.685 0.980 ;
        RECT  0.000 -0.130 0.445 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 1.890 6.845 3.000 ;
        RECT  4.795 2.740 6.585 3.000 ;
        RECT  4.535 2.305 4.795 3.000 ;
        RECT  2.105 2.740 4.535 3.000 ;
        RECT  1.845 2.620 2.105 3.000 ;
        RECT  0.345 2.740 1.845 3.000 ;
        RECT  0.145 1.795 0.345 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.915 1.355 5.455 1.515 ;
        RECT  3.755 0.835 3.915 1.515 ;
        RECT  3.090 0.835 3.755 0.995 ;
        RECT  2.930 0.835 3.090 2.075 ;
        RECT  2.605 0.835 2.930 0.995 ;
        RECT  2.715 1.815 2.930 2.075 ;
        RECT  2.445 0.395 2.605 0.995 ;
        RECT  1.025 0.540 2.445 0.700 ;
        RECT  1.025 1.840 1.250 2.100 ;
        RECT  0.865 0.540 1.025 2.100 ;
    END
END OR2X12MTH

MACRO OR2X1MTH
    CLASS CORE ;
    FOREIGN OR2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.720 1.950 2.135 ;
        RECT  1.715 0.720 1.740 0.980 ;
        RECT  1.685 1.875 1.740 2.135 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.375 1.130 1.990 ;
        END
        AntennaGateArea 0.0741 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.225 0.380 1.485 ;
        RECT  0.100 0.880 0.310 1.580 ;
        END
        AntennaGateArea 0.0741 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.755 -0.130 2.050 0.130 ;
        RECT  1.415 -0.130 1.755 0.320 ;
        RECT  1.155 -0.130 1.415 1.025 ;
        RECT  0.365 -0.130 1.155 0.130 ;
        RECT  0.145 -0.130 0.365 0.690 ;
        RECT  0.000 -0.130 0.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.355 2.740 2.050 3.000 ;
        RECT  0.415 2.510 1.355 3.000 ;
        RECT  0.000 2.740 0.415 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.470 1.315 1.560 1.575 ;
        RECT  1.310 1.315 1.470 2.330 ;
        RECT  0.720 2.170 1.310 2.330 ;
        RECT  0.720 0.375 0.895 0.535 ;
        RECT  0.560 0.375 0.720 2.330 ;
        RECT  0.175 1.815 0.560 2.075 ;
    END
END OR2X1MTH

MACRO OR2X2MTH
    CLASS CORE ;
    FOREIGN OR2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.050 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 0.355 1.950 2.395 ;
        RECT  1.665 0.355 1.740 0.955 ;
        RECT  1.635 1.795 1.740 2.395 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.880 1.315 1.130 1.990 ;
        END
        AntennaGateArea 0.1209 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.940 0.355 1.580 ;
        END
        AntennaGateArea 0.1209 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.385 -0.130 2.050 0.130 ;
        RECT  0.785 -0.130 1.385 0.475 ;
        RECT  0.385 -0.130 0.785 0.130 ;
        RECT  0.125 -0.130 0.385 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.295 2.740 2.050 3.000 ;
        RECT  1.035 2.190 1.295 3.000 ;
        RECT  0.780 2.740 1.035 3.000 ;
        RECT  0.180 2.570 0.780 3.000 ;
        RECT  0.000 2.740 0.180 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.485 1.315 1.560 1.575 ;
        RECT  1.325 0.975 1.485 1.575 ;
        RECT  0.895 0.975 1.325 1.135 ;
        RECT  0.695 0.765 0.895 1.135 ;
        RECT  0.535 0.765 0.695 2.110 ;
        RECT  0.125 1.850 0.535 2.110 ;
    END
END OR2X2MTH

MACRO OR2X4MTH
    CLASS CORE ;
    FOREIGN OR2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.785 0.765 1.950 2.060 ;
        RECT  1.775 0.765 1.785 2.395 ;
        RECT  1.740 0.375 1.775 2.395 ;
        RECT  1.615 0.375 1.740 0.975 ;
        RECT  1.525 1.795 1.740 2.395 ;
        END
        AntennaDiffArea 0.604 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.085 1.700 1.130 1.990 ;
        RECT  0.875 1.305 1.085 1.990 ;
        END
        AntennaGateArea 0.1924 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.225 0.355 1.485 ;
        RECT  0.100 0.905 0.310 1.580 ;
        END
        AntennaGateArea 0.1924 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.335 -0.130 2.460 0.130 ;
        RECT  2.075 -0.130 2.335 0.625 ;
        RECT  0.000 -0.130 2.075 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 2.740 2.460 3.000 ;
        RECT  2.065 2.220 2.325 3.000 ;
        RECT  1.245 2.740 2.065 3.000 ;
        RECT  0.985 2.190 1.245 3.000 ;
        RECT  0.000 2.740 0.985 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.435 1.315 1.560 1.575 ;
        RECT  1.275 0.965 1.435 1.575 ;
        RECT  0.895 0.965 1.275 1.125 ;
        RECT  0.695 0.700 0.895 1.125 ;
        RECT  0.535 0.700 0.695 1.965 ;
        RECT  0.385 1.765 0.535 1.965 ;
        RECT  0.125 1.765 0.385 2.365 ;
    END
END OR2X4MTH

MACRO OR2X6MTH
    CLASS CORE ;
    FOREIGN OR2X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.730 0.385 4.000 2.415 ;
        RECT  3.715 0.385 3.730 1.040 ;
        RECT  3.715 1.660 3.730 2.415 ;
        RECT  3.010 0.770 3.715 1.040 ;
        RECT  2.920 1.660 3.715 1.930 ;
        RECT  2.740 0.385 3.010 1.040 ;
        RECT  2.660 1.660 2.920 2.415 ;
        END
        AntennaDiffArea 1.137 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.060 1.225 2.220 2.310 ;
        RECT  0.760 2.150 2.060 2.310 ;
        RECT  0.515 2.150 0.760 2.360 ;
        RECT  0.355 1.225 0.515 2.360 ;
        END
        AntennaGateArea 0.3458 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 0.880 1.540 1.395 ;
        RECT  1.035 1.135 1.330 1.395 ;
        END
        AntennaGateArea 0.3458 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 -0.130 4.100 0.130 ;
        RECT  3.205 -0.130 3.465 0.590 ;
        RECT  2.445 -0.130 3.205 0.130 ;
        RECT  2.185 -0.130 2.445 0.615 ;
        RECT  1.415 -0.130 2.185 0.130 ;
        RECT  1.155 -0.130 1.415 0.615 ;
        RECT  0.385 -0.130 1.155 0.130 ;
        RECT  0.125 -0.130 0.385 0.640 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.450 2.740 4.100 3.000 ;
        RECT  3.190 2.110 3.450 3.000 ;
        RECT  2.330 2.740 3.190 3.000 ;
        RECT  2.070 2.540 2.330 3.000 ;
        RECT  0.555 2.740 2.070 3.000 ;
        RECT  0.295 2.540 0.555 3.000 ;
        RECT  0.000 2.740 0.295 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.560 1.220 3.550 1.480 ;
        RECT  2.400 0.840 2.560 1.480 ;
        RECT  1.925 0.840 2.400 1.000 ;
        RECT  1.880 0.420 1.925 1.000 ;
        RECT  1.720 0.420 1.880 1.950 ;
        RECT  1.665 0.420 1.720 0.680 ;
        RECT  0.855 1.790 1.720 1.950 ;
        RECT  0.855 0.410 0.905 0.670 ;
        RECT  0.695 0.410 0.855 1.950 ;
        RECT  0.645 0.410 0.695 0.670 ;
    END
END OR2X6MTH

MACRO OR2X8MTH
    CLASS CORE ;
    FOREIGN OR2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.890 0.745 4.065 2.030 ;
        RECT  3.885 0.350 3.890 2.030 ;
        RECT  3.725 0.350 3.885 2.465 ;
        RECT  3.540 0.350 3.725 1.085 ;
        RECT  3.535 1.690 3.725 2.465 ;
        RECT  2.895 0.745 3.540 1.085 ;
        RECT  2.805 1.690 3.535 2.030 ;
        RECT  2.565 0.385 2.895 1.085 ;
        RECT  2.455 1.690 2.805 2.465 ;
        END
        AntennaDiffArea 1.204 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.945 1.315 2.045 1.575 ;
        RECT  1.785 1.315 1.945 2.310 ;
        RECT  0.760 2.150 1.785 2.310 ;
        RECT  0.515 2.150 0.760 2.360 ;
        RECT  0.355 1.225 0.515 2.360 ;
        RECT  0.255 1.225 0.355 1.485 ;
        END
        AntennaGateArea 0.3848 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.160 1.085 1.540 1.580 ;
        END
        AntennaGateArea 0.3848 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 -0.130 4.510 0.130 ;
        RECT  4.125 -0.130 4.385 0.560 ;
        RECT  3.335 -0.130 4.125 0.130 ;
        RECT  3.075 -0.130 3.335 0.565 ;
        RECT  0.385 -0.130 3.075 0.130 ;
        RECT  0.125 -0.130 0.385 0.755 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.385 2.740 4.510 3.000 ;
        RECT  4.125 2.215 4.385 3.000 ;
        RECT  3.300 2.740 4.125 3.000 ;
        RECT  3.040 2.215 3.300 3.000 ;
        RECT  2.210 2.740 3.040 3.000 ;
        RECT  1.950 2.570 2.210 3.000 ;
        RECT  0.455 2.740 1.950 3.000 ;
        RECT  0.195 2.620 0.455 3.000 ;
        RECT  0.000 2.740 0.195 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.385 1.305 3.490 1.465 ;
        RECT  2.225 0.735 2.385 1.465 ;
        RECT  1.865 0.735 2.225 0.895 ;
        RECT  1.605 0.495 1.865 0.895 ;
        RECT  0.855 0.735 1.605 0.895 ;
        RECT  0.855 1.790 1.325 1.950 ;
        RECT  0.695 0.495 0.855 1.950 ;
    END
END OR2X8MTH

MACRO OR3X12MTH
    CLASS CORE ;
    FOREIGN OR3X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.145 0.425 10.405 2.345 ;
        RECT  9.735 0.485 10.145 2.345 ;
        RECT  8.395 0.485 9.735 1.025 ;
        RECT  8.255 1.745 9.735 2.345 ;
        RECT  8.135 0.425 8.395 1.025 ;
        END
        AntennaDiffArea 1.8 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.590 1.265 7.590 1.540 ;
        END
        AntennaGateArea 0.8034 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.155 1.265 5.155 1.540 ;
        END
        AntennaGateArea 0.8034 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.555 1.265 2.555 1.540 ;
        END
        AntennaGateArea 0.8034 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 -0.130 11.070 0.130 ;
        RECT  10.685 -0.130 10.945 0.980 ;
        RECT  9.865 -0.130 10.685 0.130 ;
        RECT  9.605 -0.130 9.865 0.300 ;
        RECT  7.840 -0.130 9.605 0.130 ;
        RECT  7.580 -0.130 7.840 0.640 ;
        RECT  6.775 -0.130 7.580 0.130 ;
        RECT  6.515 -0.130 6.775 0.640 ;
        RECT  5.675 -0.130 6.515 0.130 ;
        RECT  5.415 -0.130 5.675 0.640 ;
        RECT  4.575 -0.130 5.415 0.130 ;
        RECT  4.315 -0.130 4.575 0.640 ;
        RECT  3.475 -0.130 4.315 0.130 ;
        RECT  3.215 -0.130 3.475 0.640 ;
        RECT  3.030 -0.130 3.215 0.130 ;
        RECT  2.770 -0.130 3.030 0.640 ;
        RECT  1.970 -0.130 2.770 0.130 ;
        RECT  1.710 -0.130 1.970 0.640 ;
        RECT  0.880 -0.130 1.710 0.130 ;
        RECT  0.620 -0.130 0.880 0.640 ;
        RECT  0.400 -0.130 0.620 0.130 ;
        RECT  0.140 -0.130 0.400 0.640 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 2.740 11.070 3.000 ;
        RECT  10.685 1.890 10.945 3.000 ;
        RECT  6.095 2.740 10.685 3.000 ;
        RECT  5.835 2.210 6.095 3.000 ;
        RECT  0.000 2.740 5.835 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.175 1.255 9.455 1.515 ;
        RECT  7.940 1.255 8.175 1.415 ;
        RECT  7.780 0.845 7.940 1.415 ;
        RECT  7.320 0.845 7.780 1.045 ;
        RECT  7.305 1.870 7.565 2.470 ;
        RECT  7.060 0.710 7.320 1.045 ;
        RECT  6.615 1.870 7.305 2.030 ;
        RECT  6.225 0.845 7.060 1.045 ;
        RECT  6.355 1.870 6.615 2.470 ;
        RECT  5.575 1.870 6.355 2.030 ;
        RECT  5.965 0.710 6.225 1.045 ;
        RECT  5.120 0.845 5.965 1.045 ;
        RECT  5.315 1.870 5.575 2.470 ;
        RECT  4.535 1.870 5.315 2.030 ;
        RECT  4.860 0.710 5.120 1.045 ;
        RECT  4.795 2.215 5.055 2.475 ;
        RECT  4.025 0.845 4.860 1.045 ;
        RECT  4.015 2.315 4.795 2.475 ;
        RECT  4.275 1.870 4.535 2.130 ;
        RECT  3.495 1.870 4.275 2.030 ;
        RECT  3.765 0.710 4.025 1.045 ;
        RECT  3.755 2.215 4.015 2.475 ;
        RECT  2.520 0.845 3.765 1.045 ;
        RECT  2.975 2.315 3.755 2.475 ;
        RECT  3.235 1.870 3.495 2.130 ;
        RECT  2.715 1.815 2.975 2.475 ;
        RECT  0.645 1.815 2.715 1.975 ;
        RECT  2.260 0.710 2.520 1.045 ;
        RECT  0.355 2.215 2.460 2.475 ;
        RECT  1.425 0.845 2.260 1.045 ;
        RECT  1.165 0.710 1.425 1.045 ;
        RECT  0.355 0.845 1.165 1.045 ;
        RECT  0.155 0.845 0.355 2.475 ;
    END
END OR3X12MTH

MACRO OR3X1MTH
    CLASS CORE ;
    FOREIGN OR3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.155 0.765 2.360 2.045 ;
        RECT  2.125 0.765 2.155 1.025 ;
        RECT  2.085 1.700 2.155 2.045 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.115 1.565 1.600 ;
        END
        AntennaGateArea 0.0871 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.830 1.115 1.130 1.600 ;
        END
        AntennaGateArea 0.0871 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.625 1.580 ;
        END
        AntennaGateArea 0.0871 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.255 -0.130 2.460 0.130 ;
        RECT  1.655 -0.130 2.255 0.415 ;
        RECT  0.865 -0.130 1.655 0.130 ;
        RECT  0.265 -0.130 0.865 0.515 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.755 2.740 2.460 3.000 ;
        RECT  1.495 2.125 1.755 3.000 ;
        RECT  1.145 2.740 1.495 3.000 ;
        RECT  0.205 2.570 1.145 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.905 1.225 1.975 1.485 ;
        RECT  1.745 0.775 1.905 1.940 ;
        RECT  1.395 0.775 1.745 0.935 ;
        RECT  0.385 1.780 1.745 1.940 ;
        RECT  1.135 0.340 1.395 0.935 ;
        RECT  0.385 0.775 1.135 0.935 ;
        RECT  0.125 0.775 0.385 0.975 ;
        RECT  0.125 1.780 0.385 2.040 ;
    END
END OR3X1MTH

MACRO OR3X2MTH
    CLASS CORE ;
    FOREIGN OR3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.460 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.180 0.390 2.360 2.385 ;
        RECT  2.125 0.390 2.180 0.990 ;
        RECT  2.125 1.700 2.180 2.385 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.155 1.600 1.600 ;
        END
        AntennaGateArea 0.1404 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.755 1.155 1.130 1.600 ;
        END
        AntennaGateArea 0.1404 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.225 0.575 1.580 ;
        END
        AntennaGateArea 0.1404 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.795 -0.130 2.460 0.130 ;
        RECT  1.195 -0.130 1.795 0.475 ;
        RECT  0.785 -0.130 1.195 0.130 ;
        RECT  0.185 -0.130 0.785 0.475 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.765 2.740 2.460 3.000 ;
        RECT  1.505 2.120 1.765 3.000 ;
        RECT  0.000 2.740 1.505 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  1.945 1.265 2.000 1.525 ;
        RECT  1.785 0.815 1.945 1.940 ;
        RECT  0.125 0.815 1.785 0.975 ;
        RECT  0.385 1.780 1.785 1.940 ;
        RECT  0.125 1.780 0.385 2.380 ;
    END
END OR3X2MTH

MACRO OR3X4MTH
    CLASS CORE ;
    FOREIGN OR3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.740 1.285 4.040 1.585 ;
        RECT  3.560 0.380 3.740 2.395 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.850 1.225 2.950 1.485 ;
        RECT  2.690 0.920 2.850 1.485 ;
        RECT  0.760 0.920 2.690 1.080 ;
        RECT  0.690 0.920 0.760 1.130 ;
        RECT  0.430 0.920 0.690 1.485 ;
        END
        AntennaGateArea 0.2821 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.210 1.295 2.470 1.950 ;
        RECT  1.170 1.740 2.210 1.950 ;
        RECT  0.910 1.320 1.170 1.950 ;
        END
        AntennaGateArea 0.2821 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.390 1.260 1.990 1.540 ;
        END
        AntennaGateArea 0.2821 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.310 -0.130 4.510 0.130 ;
        RECT  4.050 -0.130 4.310 0.980 ;
        RECT  3.215 -0.130 4.050 0.130 ;
        RECT  2.955 -0.130 3.215 0.300 ;
        RECT  1.970 -0.130 2.955 0.130 ;
        RECT  1.710 -0.130 1.970 0.300 ;
        RECT  0.745 -0.130 1.710 0.130 ;
        RECT  0.145 -0.130 0.745 0.300 ;
        RECT  0.000 -0.130 0.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.310 2.740 4.510 3.000 ;
        RECT  4.050 1.795 4.310 3.000 ;
        RECT  3.230 2.740 4.050 3.000 ;
        RECT  2.970 2.470 3.230 3.000 ;
        RECT  0.480 2.740 2.970 3.000 ;
        RECT  0.220 1.685 0.480 3.000 ;
        RECT  0.000 2.740 0.220 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.220 0.580 3.380 2.290 ;
        RECT  1.050 0.580 3.220 0.740 ;
        RECT  1.820 2.130 3.220 2.290 ;
        RECT  1.560 2.130 1.820 2.390 ;
    END
END OR3X4MTH

MACRO OR3X6MTH
    CLASS CORE ;
    FOREIGN OR3X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.920 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.540 0.380 4.820 2.395 ;
        RECT  3.685 0.805 4.540 1.015 ;
        RECT  3.685 1.795 4.540 2.005 ;
        RECT  3.425 0.380 3.685 1.015 ;
        RECT  3.425 1.795 3.685 2.395 ;
        END
        AntennaDiffArea 1.137 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.650 0.920 2.810 1.485 ;
        RECT  0.760 0.920 2.650 1.080 ;
        RECT  0.595 0.920 0.760 1.130 ;
        RECT  0.335 0.920 0.595 1.485 ;
        END
        AntennaGateArea 0.2951 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.120 1.295 2.380 1.965 ;
        RECT  1.170 1.805 2.120 1.965 ;
        RECT  1.075 1.740 1.170 1.965 ;
        RECT  0.815 1.320 1.075 1.965 ;
        END
        AntennaGateArea 0.2951 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.330 1.270 1.810 1.580 ;
        END
        AntennaGateArea 0.2951 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.225 -0.130 4.920 0.130 ;
        RECT  3.965 -0.130 4.225 0.625 ;
        RECT  3.140 -0.130 3.965 0.130 ;
        RECT  2.880 -0.130 3.140 0.400 ;
        RECT  2.005 -0.130 2.880 0.130 ;
        RECT  1.745 -0.130 2.005 0.400 ;
        RECT  0.850 -0.130 1.745 0.130 ;
        RECT  0.250 -0.130 0.850 0.300 ;
        RECT  0.000 -0.130 0.250 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.225 2.740 4.920 3.000 ;
        RECT  3.965 2.185 4.225 3.000 ;
        RECT  3.105 2.740 3.965 3.000 ;
        RECT  2.845 2.490 3.105 3.000 ;
        RECT  0.385 2.740 2.845 3.000 ;
        RECT  0.125 1.800 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.150 1.225 4.315 1.485 ;
        RECT  2.990 0.580 3.150 2.310 ;
        RECT  1.205 0.580 2.990 0.740 ;
        RECT  1.465 2.150 2.990 2.310 ;
    END
END OR3X6MTH

MACRO OR3X8MTH
    CLASS CORE ;
    FOREIGN OR3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.350 0.735 6.465 2.400 ;
        RECT  6.115 0.385 6.350 2.400 ;
        RECT  6.000 0.385 6.115 1.095 ;
        RECT  5.545 1.695 6.115 2.045 ;
        RECT  5.320 0.745 6.000 1.095 ;
        RECT  5.195 1.695 5.545 2.400 ;
        RECT  4.970 0.385 5.320 1.095 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.610 1.225 4.450 1.540 ;
        END
        AntennaGateArea 0.4979 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 1.225 3.020 1.540 ;
        END
        AntennaGateArea 0.4979 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.545 1.225 1.525 1.540 ;
        END
        AntennaGateArea 0.4979 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.835 -0.130 6.970 0.130 ;
        RECT  6.625 -0.130 6.835 0.650 ;
        RECT  5.780 -0.130 6.625 0.130 ;
        RECT  5.520 -0.130 5.780 0.565 ;
        RECT  4.625 -0.130 5.520 0.130 ;
        RECT  4.365 -0.130 4.625 0.705 ;
        RECT  3.450 -0.130 4.365 0.130 ;
        RECT  3.190 -0.130 3.450 0.705 ;
        RECT  2.370 -0.130 3.190 0.130 ;
        RECT  1.730 -0.130 2.370 0.660 ;
        RECT  1.500 -0.130 1.730 0.130 ;
        RECT  1.240 -0.130 1.500 0.660 ;
        RECT  0.385 -0.130 1.240 0.130 ;
        RECT  0.125 -0.130 0.385 0.705 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.975 2.740 6.970 3.000 ;
        RECT  4.715 1.890 4.975 3.000 ;
        RECT  0.000 2.740 4.715 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.790 1.315 5.935 1.475 ;
        RECT  4.630 0.885 4.790 1.475 ;
        RECT  4.000 0.885 4.630 1.045 ;
        RECT  4.165 1.875 4.425 2.475 ;
        RECT  3.475 1.875 4.165 2.035 ;
        RECT  3.740 0.515 4.000 1.045 ;
        RECT  2.900 0.885 3.740 1.045 ;
        RECT  3.215 1.875 3.475 2.475 ;
        RECT  2.435 1.875 3.215 2.035 ;
        RECT  2.695 2.215 2.955 2.475 ;
        RECT  2.640 0.515 2.900 1.045 ;
        RECT  1.915 2.315 2.695 2.475 ;
        RECT  0.930 0.885 2.640 1.045 ;
        RECT  2.175 1.875 2.435 2.135 ;
        RECT  1.655 1.875 1.915 2.475 ;
        RECT  0.895 1.875 1.655 2.035 ;
        RECT  0.365 2.215 1.370 2.475 ;
        RECT  0.670 0.640 0.930 1.045 ;
        RECT  0.635 1.775 0.895 2.035 ;
        RECT  0.365 0.885 0.670 1.045 ;
        RECT  0.145 0.885 0.365 2.475 ;
    END
END OR3X8MTH

MACRO OR4X12MTH
    CLASS CORE ;
    FOREIGN OR4X12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.450 0.380 13.710 2.345 ;
        RECT  13.015 0.745 13.450 2.125 ;
        RECT  12.690 0.745 13.015 1.135 ;
        RECT  12.690 1.735 13.015 2.125 ;
        RECT  12.430 0.380 12.690 1.135 ;
        RECT  12.430 1.735 12.690 2.345 ;
        RECT  11.710 0.745 12.430 1.135 ;
        RECT  11.670 1.735 12.430 2.125 ;
        RECT  11.450 0.405 11.710 1.135 ;
        RECT  11.410 1.735 11.670 2.345 ;
        RECT  10.690 0.745 11.450 1.135 ;
        RECT  10.430 0.405 10.690 1.135 ;
        END
        AntennaDiffArea 1.865 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.215 2.035 1.475 ;
        RECT  0.920 1.215 1.130 1.580 ;
        RECT  0.515 1.215 0.920 1.475 ;
        END
        AntennaGateArea 0.8502 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.225 4.680 1.485 ;
        RECT  4.200 1.225 4.410 1.580 ;
        RECT  3.160 1.225 4.200 1.485 ;
        END
        AntennaGateArea 0.8502 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.870 1.225 7.850 1.485 ;
        RECT  6.660 1.225 6.870 1.580 ;
        RECT  6.330 1.225 6.660 1.485 ;
        END
        AntennaGateArea 0.8502 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.920 1.225 9.860 1.485 ;
        RECT  8.710 1.225 8.920 1.580 ;
        RECT  8.340 1.225 8.710 1.485 ;
        END
        AntennaGateArea 0.8502 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.220 -0.130 14.350 0.130 ;
        RECT  13.960 -0.130 14.220 0.970 ;
        RECT  13.200 -0.130 13.960 0.130 ;
        RECT  12.940 -0.130 13.200 0.565 ;
        RECT  11.200 -0.130 12.940 0.130 ;
        RECT  10.940 -0.130 11.200 0.565 ;
        RECT  6.830 -0.130 10.940 0.130 ;
        RECT  6.570 -0.130 6.830 0.565 ;
        RECT  6.235 -0.130 6.570 0.130 ;
        RECT  5.635 -0.130 6.235 0.300 ;
        RECT  5.315 -0.130 5.635 0.130 ;
        RECT  5.055 -0.130 5.315 0.605 ;
        RECT  1.425 -0.130 5.055 0.130 ;
        RECT  1.165 -0.130 1.425 0.615 ;
        RECT  0.385 -0.130 1.165 0.130 ;
        RECT  0.125 -0.130 0.385 0.745 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.220 2.740 14.350 3.000 ;
        RECT  13.960 1.865 14.220 3.000 ;
        RECT  13.200 2.740 13.960 3.000 ;
        RECT  12.940 2.305 13.200 3.000 ;
        RECT  12.180 2.740 12.940 3.000 ;
        RECT  11.920 2.305 12.180 3.000 ;
        RECT  11.160 2.740 11.920 3.000 ;
        RECT  10.900 2.255 11.160 3.000 ;
        RECT  2.465 2.740 10.900 3.000 ;
        RECT  2.205 2.255 2.465 3.000 ;
        RECT  1.425 2.740 2.205 3.000 ;
        RECT  1.165 2.255 1.425 3.000 ;
        RECT  0.385 2.740 1.165 3.000 ;
        RECT  0.125 1.850 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.030 1.355 12.730 1.515 ;
        RECT  10.770 1.355 11.030 1.945 ;
        RECT  10.220 1.685 10.770 1.945 ;
        RECT  9.990 2.215 10.250 2.475 ;
        RECT  10.180 0.785 10.220 1.945 ;
        RECT  10.060 0.365 10.180 1.945 ;
        RECT  9.920 0.365 10.060 0.955 ;
        RECT  9.740 1.785 10.060 1.945 ;
        RECT  9.230 2.315 9.990 2.475 ;
        RECT  9.230 0.795 9.920 0.955 ;
        RECT  9.480 1.785 9.740 2.045 ;
        RECT  8.720 1.785 9.480 1.945 ;
        RECT  8.970 0.355 9.230 0.955 ;
        RECT  8.970 2.215 9.230 2.475 ;
        RECT  8.300 0.795 8.970 0.955 ;
        RECT  8.210 2.315 8.970 2.475 ;
        RECT  8.460 1.785 8.720 2.045 ;
        RECT  8.040 0.545 8.300 0.955 ;
        RECT  7.950 1.875 8.210 2.475 ;
        RECT  7.350 0.795 8.040 0.955 ;
        RECT  7.170 2.315 7.950 2.475 ;
        RECT  7.430 1.875 7.690 2.135 ;
        RECT  6.650 1.875 7.430 2.035 ;
        RECT  7.090 0.545 7.350 0.955 ;
        RECT  6.910 2.215 7.170 2.475 ;
        RECT  4.795 0.795 7.090 0.955 ;
        RECT  6.110 2.315 6.910 2.475 ;
        RECT  6.390 1.875 6.650 2.135 ;
        RECT  5.590 1.875 6.390 2.035 ;
        RECT  5.850 2.215 6.110 2.475 ;
        RECT  5.330 1.875 5.590 2.135 ;
        RECT  4.550 1.875 5.330 2.035 ;
        RECT  4.810 2.215 5.070 2.475 ;
        RECT  4.030 2.315 4.810 2.475 ;
        RECT  4.535 0.395 4.795 0.955 ;
        RECT  4.290 1.875 4.550 2.135 ;
        RECT  3.845 0.795 4.535 0.955 ;
        RECT  3.510 1.875 4.290 2.035 ;
        RECT  3.770 2.215 4.030 2.475 ;
        RECT  3.585 0.395 3.845 0.955 ;
        RECT  2.985 2.315 3.770 2.475 ;
        RECT  2.895 0.795 3.585 0.955 ;
        RECT  3.250 1.875 3.510 2.135 ;
        RECT  2.725 1.875 2.985 2.475 ;
        RECT  2.635 0.395 2.895 0.955 ;
        RECT  1.945 1.875 2.725 2.035 ;
        RECT  1.945 0.795 2.635 0.955 ;
        RECT  1.685 0.395 1.945 0.955 ;
        RECT  1.685 1.875 1.945 2.475 ;
        RECT  0.905 0.795 1.685 0.955 ;
        RECT  0.905 1.875 1.685 2.035 ;
        RECT  0.645 0.545 0.905 0.955 ;
        RECT  0.645 1.875 0.905 2.475 ;
    END
END OR4X12MTH

MACRO OR4X1MTH
    CLASS CORE ;
    FOREIGN OR4X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.870 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.695 1.700 2.770 2.120 ;
        RECT  2.535 0.735 2.695 2.120 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.585 1.185 1.950 1.735 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.605 1.370 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.220 0.925 1.380 ;
        RECT  0.100 0.880 0.310 1.380 ;
        END
        AntennaGateArea 0.0884 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.195 1.605 0.720 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.615 -0.130 2.870 0.130 ;
        RECT  2.015 -0.130 2.615 0.300 ;
        RECT  1.255 -0.130 2.015 0.130 ;
        RECT  0.655 -0.130 1.255 0.300 ;
        RECT  0.385 -0.130 0.655 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.400 2.740 2.870 3.000 ;
        RECT  1.800 2.570 2.400 3.000 ;
        RECT  0.000 2.740 1.800 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.165 0.835 2.325 2.330 ;
        RECT  1.765 0.835 2.165 0.995 ;
        RECT  0.135 2.170 2.165 2.330 ;
        RECT  1.505 0.315 1.765 0.995 ;
        RECT  0.815 0.835 1.505 0.995 ;
        RECT  0.555 0.735 0.815 0.995 ;
    END
END OR4X1MTH

MACRO OR4X2MTH
    CLASS CORE ;
    FOREIGN OR4X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.280 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.040 0.760 3.180 2.400 ;
        RECT  2.970 0.370 3.040 2.400 ;
        RECT  2.880 0.370 2.970 0.970 ;
        RECT  2.605 2.110 2.970 2.400 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.225 2.360 1.585 ;
        END
        AntennaGateArea 0.1417 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.180 1.695 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.105 1.700 1.130 1.990 ;
        RECT  0.945 1.160 1.105 1.990 ;
        RECT  0.920 1.700 0.945 1.990 ;
        END
        AntennaGateArea 0.1417 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.225 0.620 1.545 ;
        RECT  0.100 0.880 0.310 1.545 ;
        END
        AntennaGateArea 0.1417 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.550 -0.130 3.280 0.130 ;
        RECT  1.950 -0.130 2.550 0.300 ;
        RECT  1.595 -0.130 1.950 0.130 ;
        RECT  0.995 -0.130 1.595 0.300 ;
        RECT  0.725 -0.130 0.995 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.325 2.740 3.280 3.000 ;
        RECT  2.065 2.190 2.325 3.000 ;
        RECT  0.000 2.740 2.065 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.540 0.815 2.700 1.925 ;
        RECT  0.645 0.815 2.540 0.975 ;
        RECT  1.840 1.765 2.540 1.925 ;
        RECT  1.680 1.765 1.840 2.405 ;
        RECT  0.500 2.245 1.680 2.405 ;
        RECT  0.240 1.805 0.500 2.405 ;
    END
END OR4X2MTH

MACRO OR4X4MTH
    CLASS CORE ;
    FOREIGN OR4X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.990 1.290 6.050 1.580 ;
        RECT  5.855 0.785 5.990 2.415 ;
        RECT  5.810 0.365 5.855 2.415 ;
        RECT  5.675 0.365 5.810 0.965 ;
        RECT  5.685 1.815 5.810 2.415 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.225 1.110 1.485 ;
        RECT  0.510 1.225 0.720 1.580 ;
        END
        AntennaGateArea 0.2873 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.945 1.290 2.375 1.590 ;
        END
        AntennaGateArea 0.2873 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.290 3.120 1.580 ;
        END
        AntennaGateArea 0.2873 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.210 4.480 1.500 ;
        RECT  4.200 1.210 4.410 1.580 ;
        RECT  3.980 1.210 4.200 1.500 ;
        END
        AntennaGateArea 0.2873 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.980 ;
        RECT  5.305 -0.130 6.175 0.130 ;
        RECT  5.145 -0.130 5.305 0.980 ;
        RECT  4.840 -0.130 5.145 0.130 ;
        RECT  4.240 -0.130 4.840 0.300 ;
        RECT  3.410 -0.130 4.240 0.130 ;
        RECT  3.150 -0.130 3.410 0.300 ;
        RECT  2.960 -0.130 3.150 0.130 ;
        RECT  2.360 -0.130 2.960 0.300 ;
        RECT  2.175 -0.130 2.360 0.130 ;
        RECT  1.915 -0.130 2.175 0.300 ;
        RECT  1.075 -0.130 1.915 0.130 ;
        RECT  0.815 -0.130 1.075 0.980 ;
        RECT  0.135 -0.130 0.815 0.300 ;
        RECT  0.000 -0.130 0.135 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.785 6.435 3.000 ;
        RECT  5.385 2.740 6.175 3.000 ;
        RECT  5.225 1.685 5.385 3.000 ;
        RECT  5.125 1.685 5.225 1.945 ;
        RECT  0.905 2.740 5.225 3.000 ;
        RECT  0.645 2.195 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.820 1.225 5.630 1.485 ;
        RECT  4.665 2.195 4.925 2.455 ;
        RECT  4.660 0.595 4.820 2.015 ;
        RECT  3.905 2.295 4.665 2.455 ;
        RECT  3.960 0.595 4.660 0.755 ;
        RECT  4.415 1.855 4.660 2.015 ;
        RECT  4.155 1.855 4.415 2.115 ;
        RECT  3.700 0.495 3.960 0.755 ;
        RECT  3.645 2.195 3.905 2.455 ;
        RECT  1.625 0.595 3.700 0.755 ;
        RECT  2.865 2.295 3.645 2.455 ;
        RECT  3.300 0.950 3.460 2.115 ;
        RECT  1.765 0.950 3.300 1.110 ;
        RECT  3.125 1.855 3.300 2.115 ;
        RECT  2.705 1.760 2.865 2.455 ;
        RECT  2.605 1.760 2.705 1.920 ;
        RECT  2.205 2.220 2.465 2.480 ;
        RECT  1.425 2.320 2.205 2.480 ;
        RECT  1.765 1.855 1.945 2.115 ;
        RECT  1.605 0.950 1.765 2.115 ;
        RECT  1.365 0.495 1.625 0.755 ;
        RECT  1.165 1.805 1.425 2.480 ;
        RECT  0.385 1.805 1.165 1.965 ;
        RECT  0.125 1.805 0.385 2.405 ;
    END
END OR4X4MTH

MACRO OR4X6MTH
    CLASS CORE ;
    FOREIGN OR4X6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.830 0.425 8.100 2.345 ;
        RECT  7.815 0.425 7.830 1.025 ;
        RECT  7.055 1.745 7.830 2.015 ;
        RECT  7.055 0.755 7.815 1.025 ;
        RECT  6.795 0.425 7.055 1.025 ;
        RECT  6.795 1.745 7.055 2.345 ;
        END
        AntennaDiffArea 1.137 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.640 1.225 6.040 1.485 ;
        RECT  5.430 1.225 5.640 1.580 ;
        RECT  5.200 1.225 5.430 1.485 ;
        END
        AntennaGateArea 0.4316 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.225 4.575 1.485 ;
        RECT  4.200 1.225 4.410 1.580 ;
        RECT  3.735 1.225 4.200 1.485 ;
        END
        AntennaGateArea 0.4316 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.225 3.015 1.485 ;
        RECT  2.560 1.225 2.770 1.580 ;
        RECT  2.175 1.225 2.560 1.485 ;
        END
        AntennaGateArea 0.4316 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.225 1.455 1.485 ;
        RECT  0.920 1.225 1.130 1.580 ;
        RECT  0.615 1.225 0.920 1.485 ;
        END
        AntennaGateArea 0.4316 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.530 -0.130 8.200 0.130 ;
        RECT  5.930 -0.130 6.530 0.615 ;
        RECT  5.065 -0.130 5.930 0.130 ;
        RECT  4.805 -0.130 5.065 0.615 ;
        RECT  3.915 -0.130 4.805 0.130 ;
        RECT  3.295 -0.130 3.915 0.615 ;
        RECT  2.355 -0.130 3.295 0.130 ;
        RECT  1.735 -0.130 2.355 0.615 ;
        RECT  0.860 -0.130 1.735 0.130 ;
        RECT  0.260 -0.130 0.860 0.615 ;
        RECT  0.000 -0.130 0.260 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.565 2.740 8.200 3.000 ;
        RECT  7.305 2.240 7.565 3.000 ;
        RECT  5.585 2.740 7.305 3.000 ;
        RECT  5.325 2.225 5.585 3.000 ;
        RECT  0.000 2.740 5.325 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.625 1.255 7.565 1.515 ;
        RECT  6.495 1.255 6.625 1.415 ;
        RECT  6.335 0.795 6.495 1.415 ;
        RECT  5.615 0.795 6.335 0.955 ;
        RECT  5.845 1.875 6.105 2.475 ;
        RECT  5.065 1.875 5.845 2.035 ;
        RECT  5.355 0.355 5.615 0.955 ;
        RECT  4.515 0.795 5.355 0.955 ;
        RECT  4.805 1.875 5.065 2.475 ;
        RECT  4.025 1.875 4.805 2.035 ;
        RECT  4.285 2.215 4.545 2.475 ;
        RECT  4.255 0.355 4.515 0.955 ;
        RECT  3.505 2.315 4.285 2.475 ;
        RECT  2.955 0.795 4.255 0.955 ;
        RECT  3.765 1.875 4.025 2.135 ;
        RECT  3.245 1.875 3.505 2.475 ;
        RECT  2.465 1.875 3.245 2.035 ;
        RECT  2.725 2.215 2.985 2.475 ;
        RECT  2.695 0.355 2.955 0.955 ;
        RECT  1.945 2.315 2.725 2.475 ;
        RECT  1.400 0.795 2.695 0.955 ;
        RECT  2.205 1.875 2.465 2.135 ;
        RECT  1.685 1.875 1.945 2.475 ;
        RECT  0.905 1.875 1.685 2.035 ;
        RECT  1.165 2.215 1.425 2.475 ;
        RECT  1.140 0.355 1.400 0.955 ;
        RECT  0.390 2.315 1.165 2.475 ;
        RECT  0.290 0.795 1.140 0.955 ;
        RECT  0.645 1.875 0.905 2.135 ;
        RECT  0.290 1.875 0.390 2.475 ;
        RECT  0.130 0.795 0.290 2.475 ;
    END
END OR4X6MTH

MACRO OR4X8MTH
    CLASS CORE ;
    FOREIGN OR4X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.845 0.605 10.970 1.795 ;
        RECT  10.815 0.605 10.845 2.345 ;
        RECT  10.620 0.355 10.815 2.345 ;
        RECT  10.555 0.355 10.620 0.955 ;
        RECT  10.585 1.565 10.620 2.345 ;
        RECT  9.885 1.565 10.585 1.915 ;
        RECT  9.735 0.605 10.555 0.955 ;
        RECT  9.625 1.565 9.885 2.345 ;
        RECT  9.475 0.355 9.735 0.955 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.225 2.055 1.485 ;
        RECT  0.920 1.225 1.130 1.580 ;
        RECT  0.535 1.225 0.920 1.485 ;
        END
        AntennaGateArea 0.5746 ;
    END D
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.180 1.125 3.735 1.285 ;
        RECT  2.970 1.125 3.180 1.580 ;
        RECT  2.455 1.125 2.970 1.285 ;
        END
        AntennaGateArea 0.5746 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.050 1.125 6.595 1.285 ;
        RECT  5.840 1.125 6.050 1.580 ;
        RECT  5.315 1.125 5.840 1.285 ;
        END
        AntennaGateArea 0.5746 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.690 1.225 8.585 1.485 ;
        RECT  7.480 1.225 7.690 1.580 ;
        RECT  7.065 1.225 7.480 1.485 ;
        END
        AntennaGateArea 0.5746 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 -0.130 11.480 0.130 ;
        RECT  11.095 -0.130 11.355 0.300 ;
        RECT  10.275 -0.130 11.095 0.130 ;
        RECT  10.015 -0.130 10.275 0.300 ;
        RECT  9.100 -0.130 10.015 0.130 ;
        RECT  8.500 -0.130 9.100 0.505 ;
        RECT  7.615 -0.130 8.500 0.130 ;
        RECT  7.355 -0.130 7.615 0.605 ;
        RECT  7.155 -0.130 7.355 0.130 ;
        RECT  6.895 -0.130 7.155 0.605 ;
        RECT  6.645 -0.130 6.895 0.130 ;
        RECT  6.385 -0.130 6.645 0.605 ;
        RECT  5.575 -0.130 6.385 0.130 ;
        RECT  4.940 -0.130 5.575 0.605 ;
        RECT  4.400 -0.130 4.940 0.130 ;
        RECT  3.800 -0.130 4.400 0.605 ;
        RECT  2.950 -0.130 3.800 0.130 ;
        RECT  2.690 -0.130 2.950 0.605 ;
        RECT  2.475 -0.130 2.690 0.130 ;
        RECT  2.215 -0.130 2.475 0.605 ;
        RECT  1.980 -0.130 2.215 0.130 ;
        RECT  1.720 -0.130 1.980 0.605 ;
        RECT  0.875 -0.130 1.720 0.130 ;
        RECT  0.615 -0.130 0.875 0.915 ;
        RECT  0.275 -0.130 0.615 0.300 ;
        RECT  0.000 -0.130 0.275 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 2.740 11.480 3.000 ;
        RECT  11.095 1.960 11.355 3.000 ;
        RECT  9.325 2.740 11.095 3.000 ;
        RECT  9.165 1.685 9.325 3.000 ;
        RECT  0.905 2.740 9.165 3.000 ;
        RECT  0.645 2.235 0.905 3.000 ;
        RECT  0.000 2.740 0.645 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.955 1.185 10.395 1.345 ;
        RECT  8.715 2.245 8.975 2.520 ;
        RECT  8.795 0.785 8.955 1.925 ;
        RECT  8.160 0.785 8.795 0.945 ;
        RECT  8.465 1.765 8.795 1.925 ;
        RECT  7.955 2.360 8.715 2.520 ;
        RECT  8.205 1.765 8.465 2.025 ;
        RECT  7.445 1.765 8.205 1.925 ;
        RECT  7.900 0.545 8.160 0.945 ;
        RECT  7.695 2.215 7.955 2.520 ;
        RECT  6.095 0.785 7.900 0.945 ;
        RECT  6.935 2.360 7.695 2.520 ;
        RECT  7.185 1.765 7.445 2.025 ;
        RECT  6.675 1.875 6.935 2.520 ;
        RECT  5.895 2.360 6.675 2.520 ;
        RECT  6.155 1.875 6.415 2.135 ;
        RECT  5.375 1.875 6.155 2.035 ;
        RECT  5.835 0.545 6.095 0.945 ;
        RECT  5.635 2.215 5.895 2.520 ;
        RECT  3.505 0.785 5.835 0.945 ;
        RECT  4.855 2.360 5.635 2.520 ;
        RECT  5.215 1.875 5.375 2.135 ;
        RECT  5.055 1.455 5.215 2.135 ;
        RECT  3.995 1.455 5.055 1.615 ;
        RECT  4.695 1.795 4.855 2.520 ;
        RECT  4.595 1.795 4.695 1.955 ;
        RECT  4.195 2.255 4.455 2.520 ;
        RECT  3.415 2.360 4.195 2.520 ;
        RECT  3.835 1.455 3.995 2.135 ;
        RECT  3.675 1.875 3.835 2.135 ;
        RECT  2.895 1.875 3.675 2.035 ;
        RECT  3.245 0.545 3.505 0.945 ;
        RECT  3.155 2.215 3.415 2.520 ;
        RECT  1.425 0.785 3.245 0.945 ;
        RECT  2.375 2.360 3.155 2.520 ;
        RECT  2.635 1.875 2.895 2.135 ;
        RECT  2.115 1.875 2.375 2.520 ;
        RECT  1.425 1.875 2.115 2.035 ;
        RECT  1.165 0.545 1.425 0.945 ;
        RECT  1.165 1.875 1.425 2.475 ;
        RECT  0.390 1.875 1.165 2.035 ;
        RECT  0.130 1.875 0.390 2.475 ;
    END
END OR4X8MTH

MACRO SDFFHQNX1MTH
    CLASS CORE ;
    FOREIGN SDFFHQNX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.190 1.300 1.450 ;
        RECT  0.900 1.140 1.250 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 2.060 2.230 2.245 ;
        RECT  1.590 2.060 1.970 2.220 ;
        RECT  1.430 1.760 1.590 2.220 ;
        RECT  0.720 1.760 1.430 1.920 ;
        RECT  0.560 1.140 0.720 1.920 ;
        RECT  0.510 1.165 0.560 1.580 ;
        RECT  0.430 1.165 0.510 1.525 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.170 0.735 11.380 2.125 ;
        RECT  11.095 0.735 11.170 0.995 ;
        RECT  11.095 1.865 11.170 2.125 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 2.105 3.220 2.390 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 1.115 4.860 1.540 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.295 -0.130 11.480 0.130 ;
        RECT  10.695 -0.130 11.295 0.350 ;
        RECT  10.010 -0.130 10.695 0.130 ;
        RECT  9.750 -0.130 10.010 0.250 ;
        RECT  8.580 -0.130 9.750 0.130 ;
        RECT  7.980 -0.130 8.580 0.250 ;
        RECT  6.840 -0.130 7.980 0.130 ;
        RECT  6.240 -0.130 6.840 0.250 ;
        RECT  3.255 -0.130 6.240 0.130 ;
        RECT  2.655 -0.130 3.255 0.250 ;
        RECT  1.510 -0.130 2.655 0.130 ;
        RECT  0.960 -0.130 1.510 0.495 ;
        RECT  0.740 -0.130 0.960 0.130 ;
        RECT  0.140 -0.130 0.740 0.495 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.325 2.740 11.480 3.000 ;
        RECT  10.725 2.620 11.325 3.000 ;
        RECT  8.315 2.740 10.725 3.000 ;
        RECT  7.375 2.620 8.315 3.000 ;
        RECT  3.195 2.740 7.375 3.000 ;
        RECT  2.255 2.570 3.195 3.000 ;
        RECT  0.910 2.740 2.255 3.000 ;
        RECT  0.310 2.570 0.910 3.000 ;
        RECT  0.000 2.740 0.310 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.335 1.255 10.920 1.515 ;
        RECT  10.325 2.285 10.585 2.475 ;
        RECT  10.255 0.395 10.515 0.590 ;
        RECT  10.335 0.770 10.385 0.930 ;
        RECT  10.175 0.770 10.335 2.105 ;
        RECT  9.995 2.315 10.325 2.475 ;
        RECT  9.935 0.430 10.255 0.590 ;
        RECT  10.125 0.770 10.175 0.930 ;
        RECT  9.935 1.210 9.995 2.475 ;
        RECT  9.835 0.430 9.935 2.475 ;
        RECT  9.775 0.430 9.835 1.370 ;
        RECT  9.305 2.000 9.835 2.210 ;
        RECT  9.475 0.430 9.775 0.590 ;
        RECT  9.495 1.520 9.655 1.780 ;
        RECT  9.195 1.520 9.495 1.680 ;
        RECT  9.215 0.355 9.475 0.590 ;
        RECT  9.145 1.950 9.305 2.210 ;
        RECT  9.035 1.475 9.195 1.680 ;
        RECT  9.030 1.475 9.035 1.635 ;
        RECT  8.870 0.430 9.030 1.635 ;
        RECT  8.965 2.370 9.015 2.530 ;
        RECT  8.755 2.280 8.965 2.530 ;
        RECT  7.550 0.430 8.870 0.590 ;
        RECT  8.655 1.475 8.870 1.635 ;
        RECT  7.105 2.280 8.755 2.440 ;
        RECT  8.265 1.940 8.745 2.100 ;
        RECT  8.265 0.785 8.690 0.945 ;
        RECT  8.495 1.425 8.655 1.685 ;
        RECT  8.105 0.785 8.265 2.100 ;
        RECT  7.445 1.940 8.105 2.100 ;
        RECT  7.785 1.560 7.925 1.720 ;
        RECT  7.625 0.770 7.785 1.720 ;
        RECT  6.745 0.770 7.625 0.930 ;
        RECT  7.290 0.340 7.550 0.590 ;
        RECT  7.285 1.280 7.445 2.100 ;
        RECT  6.405 0.430 7.290 0.590 ;
        RECT  7.165 1.280 7.285 1.440 ;
        RECT  6.945 1.620 7.105 2.515 ;
        RECT  6.685 1.620 6.945 1.780 ;
        RECT  3.560 2.355 6.945 2.515 ;
        RECT  6.585 0.770 6.745 1.150 ;
        RECT  6.505 1.990 6.745 2.150 ;
        RECT  6.505 0.990 6.585 1.150 ;
        RECT  6.345 0.990 6.505 2.150 ;
        RECT  6.245 0.430 6.405 0.810 ;
        RECT  5.840 0.990 6.345 1.150 ;
        RECT  5.615 0.650 6.245 0.810 ;
        RECT  3.615 0.310 6.060 0.470 ;
        RECT  5.615 1.620 5.990 1.780 ;
        RECT  5.455 0.650 5.615 2.175 ;
        RECT  5.380 0.705 5.455 0.965 ;
        RECT  3.900 2.015 5.455 2.175 ;
        RECT  5.200 1.350 5.275 1.610 ;
        RECT  5.040 0.760 5.200 1.610 ;
        RECT  4.515 0.760 5.040 0.920 ;
        RECT  4.390 0.660 4.515 0.920 ;
        RECT  4.390 1.675 4.445 1.835 ;
        RECT  4.230 0.660 4.390 1.835 ;
        RECT  4.185 1.675 4.230 1.835 ;
        RECT  3.795 0.680 3.955 1.190 ;
        RECT  3.740 1.645 3.900 2.175 ;
        RECT  3.560 1.030 3.795 1.190 ;
        RECT  3.455 0.310 3.615 0.590 ;
        RECT  3.400 1.030 3.560 2.515 ;
        RECT  2.440 0.430 3.455 0.590 ;
        RECT  2.780 0.770 2.880 0.930 ;
        RECT  2.620 0.770 2.780 1.925 ;
        RECT  2.390 1.665 2.620 1.925 ;
        RECT  2.280 0.430 2.440 0.880 ;
        RECT  2.260 0.720 2.280 0.880 ;
        RECT  2.125 0.720 2.260 1.230 ;
        RECT  2.100 0.720 2.125 1.875 ;
        RECT  1.910 0.310 2.100 0.470 ;
        RECT  1.965 1.070 2.100 1.875 ;
        RECT  1.770 1.715 1.965 1.875 ;
        RECT  1.750 0.310 1.910 0.880 ;
        RECT  0.345 0.720 1.750 0.880 ;
        RECT  1.250 2.400 1.660 2.560 ;
        RECT  1.090 2.125 1.250 2.560 ;
        RECT  0.335 2.125 1.090 2.285 ;
        RECT  0.250 0.720 0.345 1.005 ;
        RECT  0.250 1.705 0.335 2.285 ;
        RECT  0.090 0.720 0.250 2.285 ;
    END
END SDFFHQNX1MTH

MACRO SDFFHQNX2MTH
    CLASS CORE ;
    FOREIGN SDFFHQNX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.250 1.190 1.300 1.450 ;
        RECT  0.900 1.140 1.250 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.970 2.060 2.230 2.245 ;
        RECT  1.590 2.060 1.970 2.220 ;
        RECT  1.430 1.760 1.590 2.220 ;
        RECT  0.720 1.760 1.430 1.920 ;
        RECT  0.560 1.140 0.720 1.920 ;
        RECT  0.510 1.165 0.560 1.580 ;
        RECT  0.430 1.165 0.510 1.525 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.170 0.405 11.380 2.360 ;
        RECT  11.095 0.405 11.170 1.005 ;
        RECT  11.095 1.760 11.170 2.360 ;
        END
        AntennaDiffArea 0.521 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 2.105 3.220 2.390 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.570 1.115 4.905 1.540 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.815 -0.130 11.480 0.130 ;
        RECT  10.215 -0.130 10.815 0.300 ;
        RECT  10.005 -0.130 10.215 0.130 ;
        RECT  9.745 -0.130 10.005 0.250 ;
        RECT  8.445 -0.130 9.745 0.130 ;
        RECT  7.845 -0.130 8.445 0.250 ;
        RECT  7.085 -0.130 7.845 0.130 ;
        RECT  6.485 -0.130 7.085 0.250 ;
        RECT  3.350 -0.130 6.485 0.130 ;
        RECT  2.410 -0.130 3.350 0.250 ;
        RECT  1.510 -0.130 2.410 0.130 ;
        RECT  0.960 -0.130 1.510 0.495 ;
        RECT  0.740 -0.130 0.960 0.130 ;
        RECT  0.140 -0.130 0.740 0.495 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.325 2.740 11.480 3.000 ;
        RECT  9.725 2.295 10.325 3.000 ;
        RECT  8.315 2.740 9.725 3.000 ;
        RECT  7.375 2.620 8.315 3.000 ;
        RECT  3.195 2.740 7.375 3.000 ;
        RECT  2.255 2.570 3.195 3.000 ;
        RECT  2.045 2.740 2.255 3.000 ;
        RECT  1.845 2.570 2.045 3.000 ;
        RECT  0.910 2.740 1.845 3.000 ;
        RECT  0.310 2.570 0.910 3.000 ;
        RECT  0.000 2.740 0.310 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.915 1.315 10.990 1.575 ;
        RECT  10.755 0.770 10.915 1.865 ;
        RECT  10.155 0.770 10.755 0.930 ;
        RECT  10.295 1.705 10.755 1.865 ;
        RECT  9.955 1.140 10.515 1.300 ;
        RECT  10.135 1.705 10.295 1.965 ;
        RECT  9.795 0.430 9.955 2.115 ;
        RECT  9.490 0.430 9.795 0.590 ;
        RECT  9.085 1.955 9.795 2.115 ;
        RECT  9.455 1.515 9.615 1.775 ;
        RECT  9.230 0.355 9.490 0.590 ;
        RECT  9.045 1.515 9.455 1.675 ;
        RECT  8.865 1.955 9.085 2.215 ;
        RECT  8.885 0.430 9.045 1.675 ;
        RECT  8.875 0.430 8.885 0.590 ;
        RECT  8.615 0.405 8.875 0.590 ;
        RECT  8.695 2.370 8.735 2.530 ;
        RECT  8.265 0.785 8.705 0.945 ;
        RECT  8.475 2.280 8.695 2.530 ;
        RECT  7.595 0.430 8.615 0.590 ;
        RECT  8.265 1.940 8.565 2.100 ;
        RECT  7.105 2.280 8.475 2.440 ;
        RECT  8.105 0.785 8.265 2.100 ;
        RECT  7.445 1.940 8.105 2.100 ;
        RECT  7.785 1.560 7.925 1.720 ;
        RECT  7.625 0.770 7.785 1.720 ;
        RECT  6.985 0.770 7.625 0.930 ;
        RECT  7.335 0.340 7.595 0.590 ;
        RECT  7.285 1.250 7.445 2.100 ;
        RECT  6.645 0.430 7.335 0.590 ;
        RECT  7.165 1.250 7.285 1.410 ;
        RECT  6.945 1.620 7.105 2.515 ;
        RECT  6.825 0.770 6.985 1.150 ;
        RECT  6.595 1.620 6.945 1.780 ;
        RECT  3.665 2.355 6.945 2.515 ;
        RECT  6.415 0.990 6.825 1.150 ;
        RECT  6.415 1.990 6.745 2.150 ;
        RECT  6.485 0.430 6.645 0.810 ;
        RECT  5.705 0.650 6.485 0.810 ;
        RECT  6.255 0.990 6.415 2.150 ;
        RECT  3.710 0.310 6.305 0.470 ;
        RECT  5.885 0.990 6.255 1.150 ;
        RECT  5.705 1.620 6.025 1.780 ;
        RECT  5.545 0.650 5.705 2.175 ;
        RECT  5.425 0.705 5.545 0.965 ;
        RECT  4.005 2.015 5.545 2.175 ;
        RECT  5.245 1.350 5.350 1.610 ;
        RECT  5.085 0.760 5.245 1.610 ;
        RECT  4.635 0.760 5.085 0.920 ;
        RECT  4.390 0.660 4.635 0.920 ;
        RECT  4.390 1.675 4.445 1.835 ;
        RECT  4.230 0.660 4.390 1.835 ;
        RECT  4.185 1.675 4.230 1.835 ;
        RECT  3.890 0.680 4.050 1.190 ;
        RECT  3.845 1.425 4.005 2.175 ;
        RECT  3.665 1.030 3.890 1.190 ;
        RECT  3.550 0.310 3.710 0.590 ;
        RECT  3.505 1.030 3.665 2.515 ;
        RECT  2.440 0.430 3.550 0.590 ;
        RECT  2.780 0.770 2.880 0.930 ;
        RECT  2.620 0.770 2.780 1.925 ;
        RECT  2.390 1.665 2.620 1.925 ;
        RECT  2.280 0.430 2.440 0.880 ;
        RECT  2.260 0.720 2.280 0.880 ;
        RECT  2.125 0.720 2.260 1.230 ;
        RECT  2.100 0.720 2.125 1.875 ;
        RECT  1.910 0.310 2.100 0.470 ;
        RECT  1.965 1.070 2.100 1.875 ;
        RECT  1.770 1.715 1.965 1.875 ;
        RECT  1.750 0.310 1.910 0.880 ;
        RECT  0.345 0.720 1.750 0.880 ;
        RECT  1.250 2.400 1.660 2.560 ;
        RECT  1.090 2.125 1.250 2.560 ;
        RECT  0.335 2.125 1.090 2.285 ;
        RECT  0.250 0.720 0.345 1.005 ;
        RECT  0.250 1.705 0.335 2.285 ;
        RECT  0.090 0.720 0.250 2.285 ;
    END
END SDFFHQNX2MTH

MACRO SDFFHQNX4MTH
    CLASS CORE ;
    FOREIGN SDFFHQNX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 1.140 1.250 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.730 2.060 1.990 2.245 ;
        RECT  1.350 2.060 1.730 2.220 ;
        RECT  1.190 1.760 1.350 2.220 ;
        RECT  0.720 1.760 1.190 1.920 ;
        RECT  0.560 1.140 0.720 1.920 ;
        RECT  0.510 1.165 0.560 1.580 ;
        RECT  0.430 1.165 0.510 1.525 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.250 1.240 11.380 1.580 ;
        RECT  11.040 0.405 11.250 2.360 ;
        RECT  10.965 0.405 11.040 1.005 ;
        RECT  10.965 1.760 11.040 2.360 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.190 2.105 2.810 2.390 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.145 4.450 1.540 ;
        RECT  4.120 1.145 4.160 1.505 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 -0.130 11.890 0.130 ;
        RECT  11.505 -0.130 11.765 0.990 ;
        RECT  10.685 -0.130 11.505 0.130 ;
        RECT  10.425 -0.130 10.685 0.640 ;
        RECT  9.945 -0.130 10.425 0.130 ;
        RECT  9.345 -0.130 9.945 0.250 ;
        RECT  7.940 -0.130 9.345 0.130 ;
        RECT  7.340 -0.130 7.940 0.250 ;
        RECT  6.430 -0.130 7.340 0.130 ;
        RECT  5.830 -0.130 6.430 0.250 ;
        RECT  2.925 -0.130 5.830 0.130 ;
        RECT  2.325 -0.130 2.925 0.250 ;
        RECT  1.055 -0.130 2.325 0.130 ;
        RECT  0.455 -0.130 1.055 0.495 ;
        RECT  0.000 -0.130 0.455 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.765 2.740 11.890 3.000 ;
        RECT  11.505 1.775 11.765 3.000 ;
        RECT  10.685 2.740 11.505 3.000 ;
        RECT  10.425 2.175 10.685 3.000 ;
        RECT  9.460 2.740 10.425 3.000 ;
        RECT  9.260 2.395 9.460 3.000 ;
        RECT  7.545 2.740 9.260 3.000 ;
        RECT  6.945 2.620 7.545 3.000 ;
        RECT  2.790 2.740 6.945 3.000 ;
        RECT  1.850 2.570 2.790 3.000 ;
        RECT  0.665 2.740 1.850 3.000 ;
        RECT  0.405 2.570 0.665 3.000 ;
        RECT  0.000 2.740 0.405 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.695 1.220 10.795 1.480 ;
        RECT  10.535 0.820 10.695 1.845 ;
        RECT  10.115 0.820 10.535 0.980 ;
        RECT  10.145 1.685 10.535 1.845 ;
        RECT  9.510 1.190 10.250 1.450 ;
        RECT  9.900 1.685 10.145 1.945 ;
        RECT  9.855 0.720 10.115 0.980 ;
        RECT  9.690 1.685 9.900 2.555 ;
        RECT  9.640 2.395 9.690 2.555 ;
        RECT  9.350 0.430 9.510 2.070 ;
        RECT  9.010 0.430 9.350 0.590 ;
        RECT  8.570 1.910 9.350 2.070 ;
        RECT  8.570 1.470 9.140 1.730 ;
        RECT  8.750 0.355 9.010 0.590 ;
        RECT  8.410 0.430 8.570 1.730 ;
        RECT  8.410 1.910 8.570 2.210 ;
        RECT  8.400 0.430 8.410 0.590 ;
        RECT  8.140 0.340 8.400 0.590 ;
        RECT  8.235 2.400 8.370 2.560 ;
        RECT  8.025 2.280 8.235 2.560 ;
        RECT  8.070 0.770 8.230 2.100 ;
        RECT  7.140 0.430 8.140 0.590 ;
        RECT  7.970 0.770 8.070 0.930 ;
        RECT  7.035 1.940 8.070 2.100 ;
        RECT  6.645 2.280 8.025 2.440 ;
        RECT  7.730 1.245 7.890 1.505 ;
        RECT  7.375 1.245 7.730 1.405 ;
        RECT  7.215 0.770 7.375 1.405 ;
        RECT  6.330 0.770 7.215 0.930 ;
        RECT  6.880 0.310 7.140 0.590 ;
        RECT  6.875 1.140 7.035 2.100 ;
        RECT  5.990 0.430 6.880 0.590 ;
        RECT  6.595 1.140 6.875 1.300 ;
        RECT  6.485 1.595 6.645 2.515 ;
        RECT  6.185 1.595 6.485 1.755 ;
        RECT  3.255 2.355 6.485 2.515 ;
        RECT  6.170 0.770 6.330 1.150 ;
        RECT  6.005 1.990 6.305 2.150 ;
        RECT  6.005 0.990 6.170 1.150 ;
        RECT  5.845 0.990 6.005 2.150 ;
        RECT  5.830 0.430 5.990 0.810 ;
        RECT  5.430 0.990 5.845 1.150 ;
        RECT  5.130 0.650 5.830 0.810 ;
        RECT  3.260 0.310 5.650 0.470 ;
        RECT  5.130 1.545 5.480 1.805 ;
        RECT  4.970 0.650 5.130 2.175 ;
        RECT  3.595 2.015 4.970 2.175 ;
        RECT  4.630 0.805 4.790 1.345 ;
        RECT  4.150 0.805 4.630 0.965 ;
        RECT  3.940 0.705 4.150 0.965 ;
        RECT  3.940 1.675 4.040 1.835 ;
        RECT  3.780 0.705 3.940 1.835 ;
        RECT  3.435 1.565 3.595 2.175 ;
        RECT  3.430 0.680 3.590 0.980 ;
        RECT  3.255 0.820 3.430 0.980 ;
        RECT  3.100 0.310 3.260 0.590 ;
        RECT  3.095 0.820 3.255 2.515 ;
        RECT  2.200 0.430 3.100 0.590 ;
        RECT  2.540 0.770 2.640 0.930 ;
        RECT  2.380 0.770 2.540 1.875 ;
        RECT  2.100 1.715 2.380 1.875 ;
        RECT  2.040 0.430 2.200 0.880 ;
        RECT  1.790 0.720 2.040 0.880 ;
        RECT  1.395 0.310 1.860 0.470 ;
        RECT  1.630 0.720 1.790 1.875 ;
        RECT  1.530 1.715 1.630 1.875 ;
        RECT  1.010 2.400 1.420 2.560 ;
        RECT  1.235 0.310 1.395 0.880 ;
        RECT  0.345 0.720 1.235 0.880 ;
        RECT  0.850 2.125 1.010 2.560 ;
        RECT  0.335 2.125 0.850 2.285 ;
        RECT  0.250 0.720 0.345 1.005 ;
        RECT  0.250 1.735 0.335 2.285 ;
        RECT  0.090 0.720 0.250 2.285 ;
    END
END SDFFHQNX4MTH

MACRO SDFFHQNX8MTH
    CLASS CORE ;
    FOREIGN SDFFHQNX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.900 1.140 1.250 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 2.060 2.000 2.365 ;
        RECT  1.350 2.060 1.740 2.220 ;
        RECT  1.190 1.760 1.350 2.220 ;
        RECT  0.720 1.760 1.190 1.920 ;
        RECT  0.560 1.140 0.720 1.920 ;
        RECT  0.510 1.165 0.560 1.580 ;
        RECT  0.430 1.165 0.510 1.525 ;
        END
        AntennaGateArea 0.1313 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.605 0.405 12.865 2.360 ;
        RECT  12.065 1.225 12.605 1.575 ;
        RECT  11.805 0.405 12.065 2.360 ;
        RECT  11.675 0.405 11.805 1.005 ;
        RECT  11.675 1.760 11.805 2.360 ;
        END
        AntennaDiffArea 1.2 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.190 2.105 2.810 2.390 ;
        END
        AntennaGateArea 0.0988 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.145 4.450 1.540 ;
        RECT  4.120 1.145 4.160 1.505 ;
        END
        AntennaGateArea 0.1495 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 -0.130 13.530 0.130 ;
        RECT  13.145 -0.130 13.405 0.990 ;
        RECT  11.395 -0.130 13.145 0.130 ;
        RECT  11.135 -0.130 11.395 0.640 ;
        RECT  10.315 -0.130 11.135 0.130 ;
        RECT  9.715 -0.130 10.315 0.250 ;
        RECT  9.450 -0.130 9.715 0.130 ;
        RECT  8.850 -0.130 9.450 0.300 ;
        RECT  7.245 -0.130 8.850 0.130 ;
        RECT  7.045 -0.130 7.245 0.300 ;
        RECT  2.925 -0.130 7.045 0.130 ;
        RECT  2.325 -0.130 2.925 0.250 ;
        RECT  1.055 -0.130 2.325 0.130 ;
        RECT  0.455 -0.130 1.055 0.495 ;
        RECT  0.000 -0.130 0.455 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.775 13.405 3.000 ;
        RECT  11.395 2.740 13.145 3.000 ;
        RECT  10.795 2.570 11.395 3.000 ;
        RECT  10.370 2.740 10.795 3.000 ;
        RECT  10.110 1.940 10.370 3.000 ;
        RECT  9.770 2.550 10.110 3.000 ;
        RECT  9.130 2.740 9.770 3.000 ;
        RECT  8.870 2.570 9.130 3.000 ;
        RECT  7.040 2.740 8.870 3.000 ;
        RECT  6.780 2.620 7.040 3.000 ;
        RECT  2.790 2.740 6.780 3.000 ;
        RECT  1.850 2.570 2.790 3.000 ;
        RECT  0.665 2.740 1.850 3.000 ;
        RECT  0.405 2.570 0.665 3.000 ;
        RECT  0.000 2.740 0.405 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.345 1.220 11.585 1.480 ;
        RECT  11.185 0.820 11.345 1.875 ;
        RECT  10.855 0.820 11.185 0.980 ;
        RECT  10.910 1.715 11.185 1.875 ;
        RECT  10.140 1.275 11.005 1.535 ;
        RECT  10.650 1.715 10.910 1.975 ;
        RECT  10.755 0.690 10.855 0.980 ;
        RECT  10.595 0.460 10.755 0.980 ;
        RECT  9.740 0.460 10.595 0.620 ;
        RECT  9.980 0.800 10.140 1.675 ;
        RECT  8.750 0.800 9.980 0.960 ;
        RECT  9.570 1.515 9.980 1.675 ;
        RECT  8.290 1.170 9.680 1.330 ;
        RECT  9.410 1.515 9.570 2.295 ;
        RECT  9.310 2.015 9.410 2.295 ;
        RECT  8.520 2.015 9.310 2.175 ;
        RECT  8.770 1.590 9.030 1.835 ;
        RECT  7.950 1.590 8.770 1.750 ;
        RECT  8.490 0.755 8.750 0.960 ;
        RECT  7.370 2.355 8.690 2.515 ;
        RECT  8.260 1.935 8.520 2.175 ;
        RECT  8.130 0.310 8.290 1.330 ;
        RECT  7.585 0.310 8.130 0.470 ;
        RECT  8.100 1.170 8.130 1.330 ;
        RECT  7.920 1.590 7.950 2.100 ;
        RECT  7.760 0.695 7.920 2.100 ;
        RECT  7.180 1.940 7.760 2.100 ;
        RECT  7.425 0.310 7.585 0.640 ;
        RECT  7.420 0.990 7.580 1.505 ;
        RECT  6.830 0.480 7.425 0.640 ;
        RECT  6.050 0.990 7.420 1.150 ;
        RECT  7.210 2.280 7.370 2.515 ;
        RECT  6.565 2.280 7.210 2.440 ;
        RECT  7.020 1.425 7.180 2.100 ;
        RECT  6.640 1.425 7.020 1.585 ;
        RECT  6.730 0.310 6.830 0.640 ;
        RECT  6.570 0.310 6.730 0.810 ;
        RECT  5.130 0.650 6.570 0.810 ;
        RECT  6.490 2.280 6.565 2.515 ;
        RECT  6.405 2.280 6.490 2.545 ;
        RECT  6.230 2.355 6.405 2.545 ;
        RECT  3.260 0.310 6.350 0.470 ;
        RECT  6.050 1.980 6.290 2.140 ;
        RECT  5.700 2.355 6.230 2.515 ;
        RECT  5.890 0.990 6.050 2.140 ;
        RECT  5.540 1.005 5.700 2.515 ;
        RECT  3.255 2.355 5.540 2.515 ;
        RECT  5.130 1.485 5.345 1.745 ;
        RECT  4.970 0.650 5.130 2.175 ;
        RECT  3.595 2.015 4.970 2.175 ;
        RECT  4.630 0.805 4.790 1.345 ;
        RECT  4.150 0.805 4.630 0.965 ;
        RECT  3.940 0.705 4.150 0.965 ;
        RECT  3.940 1.675 4.040 1.835 ;
        RECT  3.780 0.705 3.940 1.835 ;
        RECT  3.435 1.565 3.595 2.175 ;
        RECT  3.430 0.705 3.590 0.980 ;
        RECT  3.255 0.820 3.430 0.980 ;
        RECT  3.100 0.310 3.260 0.590 ;
        RECT  3.095 0.820 3.255 2.515 ;
        RECT  2.200 0.430 3.100 0.590 ;
        RECT  2.540 0.770 2.640 0.930 ;
        RECT  2.380 0.770 2.540 1.875 ;
        RECT  2.100 1.715 2.380 1.875 ;
        RECT  2.040 0.430 2.200 0.880 ;
        RECT  1.790 0.720 2.040 0.880 ;
        RECT  1.395 0.310 1.860 0.470 ;
        RECT  1.630 0.720 1.790 1.880 ;
        RECT  1.530 1.720 1.630 1.880 ;
        RECT  1.010 2.400 1.420 2.560 ;
        RECT  1.235 0.310 1.395 0.880 ;
        RECT  0.345 0.720 1.235 0.880 ;
        RECT  0.850 2.125 1.010 2.560 ;
        RECT  0.335 2.125 0.850 2.285 ;
        RECT  0.250 0.720 0.345 1.005 ;
        RECT  0.250 1.705 0.335 2.285 ;
        RECT  0.090 0.720 0.250 2.285 ;
    END
END SDFFHQNX8MTH

MACRO SDFFHQX1MTH
    CLASS CORE ;
    FOREIGN SDFFHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.800 1.330 6.090 1.540 ;
        RECT  5.660 1.380 5.800 1.540 ;
        RECT  5.500 1.380 5.660 1.860 ;
        RECT  4.975 1.700 5.500 1.860 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.020 4.935 1.180 ;
        RECT  4.095 1.020 4.450 1.540 ;
        RECT  3.990 1.020 4.095 1.775 ;
        RECT  3.935 1.235 3.990 1.775 ;
        END
        AntennaGateArea 0.1105 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.570 1.285 12.610 1.585 ;
        RECT  12.290 0.555 12.570 2.015 ;
        RECT  12.100 1.755 12.290 2.015 ;
        END
        AntennaDiffArea 0.367 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.060 1.330 2.650 1.625 ;
        END
        AntennaGateArea 0.1053 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.355 1.735 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.075 -0.130 12.710 0.130 ;
        RECT  11.815 -0.130 12.075 0.790 ;
        RECT  10.995 -0.130 11.815 0.130 ;
        RECT  10.395 -0.130 10.995 0.250 ;
        RECT  9.315 -0.130 10.395 0.130 ;
        RECT  9.055 -0.130 9.315 0.250 ;
        RECT  7.915 -0.130 9.055 0.130 ;
        RECT  6.975 -0.130 7.915 0.250 ;
        RECT  0.355 -0.130 6.975 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.580 2.740 12.710 3.000 ;
        RECT  11.420 1.675 11.580 3.000 ;
        RECT  8.755 2.740 11.420 3.000 ;
        RECT  7.815 2.620 8.755 3.000 ;
        RECT  7.030 2.740 7.815 3.000 ;
        RECT  6.530 2.570 7.030 3.000 ;
        RECT  2.700 2.740 6.530 3.000 ;
        RECT  2.480 2.145 2.700 3.000 ;
        RECT  0.780 2.740 2.480 3.000 ;
        RECT  0.180 2.620 0.780 3.000 ;
        RECT  0.000 2.740 0.180 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.920 2.355 12.200 2.515 ;
        RECT  11.760 1.100 11.920 2.515 ;
        RECT  11.505 1.100 11.760 1.360 ;
        RECT  11.245 0.555 11.505 1.360 ;
        RECT  11.185 1.100 11.245 1.360 ;
        RECT  10.585 2.400 11.235 2.560 ;
        RECT  10.705 0.430 10.865 1.695 ;
        RECT  10.065 0.430 10.705 0.590 ;
        RECT  10.485 1.915 10.585 2.560 ;
        RECT  10.325 0.815 10.485 2.560 ;
        RECT  9.975 0.815 10.325 0.975 ;
        RECT  10.025 1.790 10.075 2.390 ;
        RECT  9.805 0.375 10.065 0.590 ;
        RECT  9.815 1.525 10.025 2.390 ;
        RECT  9.725 1.525 9.815 1.685 ;
        RECT  8.605 0.430 9.805 0.590 ;
        RECT  9.565 0.810 9.725 1.685 ;
        RECT  9.475 1.865 9.635 2.390 ;
        RECT  9.465 0.810 9.565 0.970 ;
        RECT  9.295 1.525 9.565 1.685 ;
        RECT  7.685 2.230 9.475 2.390 ;
        RECT  9.035 1.525 9.295 2.050 ;
        RECT  8.805 1.185 9.125 1.345 ;
        RECT  8.165 1.525 9.035 1.685 ;
        RECT  8.545 0.770 8.805 1.345 ;
        RECT  8.345 0.385 8.605 0.590 ;
        RECT  7.430 0.770 8.545 0.965 ;
        RECT  6.730 0.430 8.345 0.590 ;
        RECT  7.905 1.425 8.165 1.685 ;
        RECT  7.425 2.170 7.685 2.390 ;
        RECT  7.170 0.770 7.430 1.950 ;
        RECT  6.350 2.230 7.425 2.390 ;
        RECT  6.915 0.770 7.170 1.035 ;
        RECT  6.730 1.290 6.780 1.550 ;
        RECT  6.615 0.430 6.730 1.550 ;
        RECT  6.540 0.430 6.615 1.990 ;
        RECT  6.455 0.725 6.540 1.990 ;
        RECT  6.010 1.830 6.455 1.990 ;
        RECT  6.270 0.310 6.360 0.570 ;
        RECT  6.190 2.230 6.350 2.560 ;
        RECT  6.110 0.310 6.270 1.150 ;
        RECT  3.045 2.400 6.190 2.560 ;
        RECT  5.320 0.990 6.110 1.150 ;
        RECT  5.850 1.830 6.010 2.220 ;
        RECT  0.695 0.310 5.930 0.470 ;
        RECT  3.385 2.060 5.850 2.220 ;
        RECT  5.160 0.650 5.320 1.520 ;
        RECT  4.135 0.650 5.160 0.810 ;
        RECT  4.790 1.360 5.160 1.520 ;
        RECT  4.630 1.360 4.790 1.880 ;
        RECT  4.275 1.720 4.630 1.880 ;
        RECT  3.755 0.665 3.800 0.925 ;
        RECT  3.595 0.665 3.755 1.880 ;
        RECT  3.565 1.620 3.595 1.880 ;
        RECT  3.245 0.650 3.405 1.280 ;
        RECT  3.225 1.460 3.385 2.220 ;
        RECT  1.035 0.650 3.245 0.810 ;
        RECT  2.990 1.460 3.225 1.620 ;
        RECT  2.885 1.805 3.045 2.560 ;
        RECT  2.830 0.990 2.990 1.620 ;
        RECT  1.665 1.805 2.885 1.965 ;
        RECT  1.850 0.990 2.830 1.150 ;
        RECT  1.920 2.145 2.180 2.465 ;
        RECT  1.035 2.305 1.920 2.465 ;
        RECT  1.690 0.990 1.850 1.625 ;
        RECT  1.590 1.415 1.690 1.625 ;
        RECT  1.405 1.805 1.665 2.120 ;
        RECT  1.375 0.990 1.405 1.250 ;
        RECT  1.375 1.805 1.405 1.965 ;
        RECT  1.215 0.990 1.375 1.965 ;
        RECT  0.875 0.650 1.035 2.465 ;
        RECT  0.535 0.310 0.695 2.075 ;
        RECT  0.125 0.765 0.535 1.025 ;
        RECT  0.385 1.915 0.535 2.075 ;
        RECT  0.125 1.915 0.385 2.175 ;
    END
END SDFFHQX1MTH

MACRO SDFFHQX2MTH
    CLASS CORE ;
    FOREIGN SDFFHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.120 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.800 1.330 6.090 1.540 ;
        RECT  5.735 1.380 5.800 1.540 ;
        RECT  5.575 1.380 5.735 1.875 ;
        RECT  4.970 1.715 5.575 1.875 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.025 5.050 1.185 ;
        RECT  4.000 1.025 4.450 1.540 ;
        END
        AntennaGateArea 0.1261 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.735 0.405 13.000 1.540 ;
        RECT  12.435 1.260 12.735 1.540 ;
        RECT  12.275 1.260 12.435 1.985 ;
        END
        AntennaDiffArea 0.407 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.565 1.620 ;
        END
        AntennaGateArea 0.0897 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.355 1.730 ;
        END
        AntennaGateArea 0.1417 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.485 -0.130 13.120 0.130 ;
        RECT  12.225 -0.130 12.485 1.005 ;
        RECT  11.915 -0.130 12.225 0.130 ;
        RECT  11.655 -0.130 11.915 0.360 ;
        RECT  11.355 -0.130 11.655 0.130 ;
        RECT  11.195 -0.130 11.355 1.000 ;
        RECT  9.385 -0.130 11.195 0.130 ;
        RECT  9.125 -0.130 9.385 0.250 ;
        RECT  8.335 -0.130 9.125 0.130 ;
        RECT  7.735 -0.130 8.335 0.250 ;
        RECT  5.735 -0.130 7.735 0.130 ;
        RECT  5.575 -0.130 5.735 0.810 ;
        RECT  0.395 -0.130 5.575 0.130 ;
        RECT  0.235 -0.130 0.395 0.300 ;
        RECT  0.000 -0.130 0.235 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.995 2.740 13.120 3.000 ;
        RECT  12.735 1.735 12.995 3.000 ;
        RECT  11.755 2.740 12.735 3.000 ;
        RECT  11.595 1.705 11.755 3.000 ;
        RECT  8.255 2.740 11.595 3.000 ;
        RECT  7.995 2.620 8.255 3.000 ;
        RECT  7.220 2.740 7.995 3.000 ;
        RECT  6.620 2.620 7.220 3.000 ;
        RECT  2.695 2.740 6.620 3.000 ;
        RECT  2.535 2.150 2.695 3.000 ;
        RECT  0.765 2.740 2.535 3.000 ;
        RECT  0.165 2.570 0.765 3.000 ;
        RECT  0.000 2.740 0.165 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.095 2.355 12.455 2.515 ;
        RECT  11.935 1.265 12.095 2.515 ;
        RECT  11.915 1.265 11.935 1.525 ;
        RECT  11.655 0.765 11.915 1.525 ;
        RECT  11.355 1.265 11.655 1.525 ;
        RECT  11.125 2.160 11.385 2.560 ;
        RECT  10.805 2.160 11.125 2.320 ;
        RECT  11.015 1.465 11.065 1.725 ;
        RECT  10.855 0.435 11.015 1.725 ;
        RECT  10.805 0.435 10.855 0.595 ;
        RECT  10.545 0.310 10.805 0.595 ;
        RECT  10.675 1.910 10.805 2.320 ;
        RECT  10.515 1.080 10.675 2.320 ;
        RECT  8.705 0.435 10.545 0.595 ;
        RECT  10.435 1.080 10.515 1.240 ;
        RECT  9.955 2.160 10.515 2.320 ;
        RECT  10.275 0.820 10.435 1.240 ;
        RECT  10.135 1.530 10.295 1.980 ;
        RECT  10.175 0.820 10.275 0.980 ;
        RECT  9.825 1.530 10.135 1.690 ;
        RECT  9.795 1.870 9.955 2.320 ;
        RECT  9.825 0.805 9.925 0.965 ;
        RECT  9.665 0.805 9.825 1.690 ;
        RECT  9.525 1.870 9.795 2.030 ;
        RECT  8.795 1.530 9.665 1.690 ;
        RECT  9.320 2.385 9.615 2.545 ;
        RECT  9.180 1.190 9.485 1.350 ;
        RECT  9.160 2.230 9.320 2.545 ;
        RECT  9.020 0.820 9.180 1.350 ;
        RECT  7.875 2.230 9.160 2.390 ;
        RECT  7.745 0.820 9.020 0.980 ;
        RECT  8.535 1.530 8.795 2.050 ;
        RECT  8.445 0.435 8.705 0.640 ;
        RECT  8.185 1.530 8.535 1.700 ;
        RECT  7.435 0.435 8.445 0.595 ;
        RECT  8.025 1.195 8.185 1.700 ;
        RECT  7.925 1.195 8.025 1.355 ;
        RECT  7.615 2.230 7.875 2.480 ;
        RECT  7.585 0.820 7.745 1.950 ;
        RECT  6.440 2.230 7.615 2.390 ;
        RECT  7.095 0.820 7.585 0.980 ;
        RECT  7.295 1.690 7.585 1.950 ;
        RECT  7.275 0.380 7.435 0.595 ;
        RECT  6.755 0.380 7.275 0.540 ;
        RECT  6.935 0.720 7.095 0.980 ;
        RECT  6.755 1.290 6.805 1.550 ;
        RECT  6.595 0.380 6.755 1.990 ;
        RECT  6.255 0.750 6.595 1.010 ;
        RECT  6.080 1.830 6.595 1.990 ;
        RECT  6.260 2.230 6.440 2.560 ;
        RECT  6.255 0.310 6.415 0.570 ;
        RECT  3.035 2.400 6.260 2.560 ;
        RECT  6.075 0.410 6.255 0.570 ;
        RECT  5.920 1.830 6.080 2.220 ;
        RECT  5.915 0.410 6.075 1.150 ;
        RECT  3.375 2.060 5.920 2.220 ;
        RECT  5.395 0.990 5.915 1.150 ;
        RECT  5.235 0.650 5.395 1.535 ;
        RECT  4.590 0.650 5.235 0.810 ;
        RECT  4.790 1.375 5.235 1.535 ;
        RECT  4.630 1.375 4.790 1.880 ;
        RECT  4.065 1.720 4.630 1.880 ;
        RECT  0.735 0.310 4.485 0.470 ;
        RECT  3.660 0.650 3.820 1.880 ;
        RECT  3.435 0.650 3.660 0.810 ;
        RECT  3.555 1.720 3.660 1.880 ;
        RECT  3.255 0.990 3.480 1.255 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.095 0.650 3.255 1.255 ;
        RECT  2.915 1.465 3.215 1.625 ;
        RECT  1.075 0.650 3.095 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.755 0.990 2.915 1.625 ;
        RECT  1.665 1.805 2.875 1.965 ;
        RECT  1.775 0.990 2.755 1.150 ;
        RECT  1.915 2.145 2.175 2.465 ;
        RECT  1.075 2.305 1.915 2.465 ;
        RECT  1.615 0.990 1.775 1.625 ;
        RECT  1.415 1.805 1.665 2.120 ;
        RECT  1.405 0.990 1.415 2.120 ;
        RECT  1.255 0.990 1.405 1.965 ;
        RECT  0.915 0.650 1.075 2.465 ;
        RECT  0.575 0.310 0.735 2.070 ;
        RECT  0.125 0.765 0.575 1.025 ;
        RECT  0.385 1.910 0.575 2.070 ;
        RECT  0.125 1.910 0.385 2.170 ;
    END
END SDFFHQX2MTH

MACRO SDFFHQX4MTH
    CLASS CORE ;
    FOREIGN SDFFHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.285 1.270 5.680 1.540 ;
        RECT  4.760 1.380 5.285 1.540 ;
        END
        AntennaGateArea 0.0806 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.035 5.070 1.195 ;
        RECT  4.220 1.035 4.450 1.540 ;
        RECT  4.060 1.035 4.220 1.725 ;
        END
        AntennaGateArea 0.1768 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.895 1.290 13.020 1.580 ;
        RECT  12.635 0.400 12.895 2.380 ;
        END
        AntennaDiffArea 0.582 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.405 1.330 2.855 1.620 ;
        END
        AntennaGateArea 0.143 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.655 1.580 ;
        END
        AntennaGateArea 0.2158 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 -0.130 13.530 0.130 ;
        RECT  13.145 -0.130 13.405 1.000 ;
        RECT  12.385 -0.130 13.145 0.130 ;
        RECT  12.125 -0.130 12.385 1.000 ;
        RECT  11.665 -0.130 12.125 0.130 ;
        RECT  11.065 -0.130 11.665 0.250 ;
        RECT  9.340 -0.130 11.065 0.130 ;
        RECT  9.080 -0.130 9.340 0.250 ;
        RECT  8.145 -0.130 9.080 0.130 ;
        RECT  7.885 -0.130 8.145 0.250 ;
        RECT  0.655 -0.130 7.885 0.130 ;
        RECT  0.495 -0.130 0.655 0.300 ;
        RECT  0.000 -0.130 0.495 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.785 13.405 3.000 ;
        RECT  12.295 2.740 13.145 3.000 ;
        RECT  11.695 2.415 12.295 3.000 ;
        RECT  9.415 2.740 11.695 3.000 ;
        RECT  9.155 2.620 9.415 3.000 ;
        RECT  8.330 2.740 9.155 3.000 ;
        RECT  8.070 2.620 8.330 3.000 ;
        RECT  2.805 2.740 8.070 3.000 ;
        RECT  2.645 2.245 2.805 3.000 ;
        RECT  2.175 2.740 2.645 3.000 ;
        RECT  1.915 2.620 2.175 3.000 ;
        RECT  0.815 2.740 1.915 3.000 ;
        RECT  0.215 2.310 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.340 1.210 12.390 1.470 ;
        RECT  12.180 1.210 12.340 2.235 ;
        RECT  12.130 1.210 12.180 1.470 ;
        RECT  10.975 2.075 12.180 2.235 ;
        RECT  11.815 1.735 11.925 1.895 ;
        RECT  11.555 0.760 11.815 1.895 ;
        RECT  11.455 1.295 11.555 1.575 ;
        RECT  11.185 1.575 11.235 1.735 ;
        RECT  11.025 0.430 11.185 1.735 ;
        RECT  10.680 0.430 11.025 0.590 ;
        RECT  10.975 1.575 11.025 1.735 ;
        RECT  10.725 1.945 10.975 2.445 ;
        RECT  10.565 0.780 10.725 2.445 ;
        RECT  10.420 0.310 10.680 0.590 ;
        RECT  10.160 0.780 10.565 0.940 ;
        RECT  9.645 2.285 10.565 2.445 ;
        RECT  6.855 0.430 10.420 0.590 ;
        RECT  10.225 1.560 10.385 1.995 ;
        RECT  9.860 1.560 10.225 1.720 ;
        RECT  9.860 0.775 9.910 0.935 ;
        RECT  9.700 0.775 9.860 1.720 ;
        RECT  9.650 0.775 9.700 0.935 ;
        RECT  8.875 1.560 9.700 1.720 ;
        RECT  9.465 1.900 9.645 2.060 ;
        RECT  9.275 1.900 9.465 2.390 ;
        RECT  7.890 2.230 9.275 2.390 ;
        RECT  9.045 1.220 9.080 1.380 ;
        RECT  8.970 1.150 9.045 1.380 ;
        RECT  8.760 0.815 8.970 1.380 ;
        RECT  8.615 1.560 8.875 2.050 ;
        RECT  7.245 0.815 8.760 0.975 ;
        RECT  8.255 1.560 8.615 1.720 ;
        RECT  7.995 1.185 8.255 1.720 ;
        RECT  7.730 2.230 7.890 2.560 ;
        RECT  3.145 2.400 7.730 2.560 ;
        RECT  7.315 1.770 7.575 2.030 ;
        RECT  7.245 1.770 7.315 1.930 ;
        RECT  7.085 0.815 7.245 1.930 ;
        RECT  7.035 0.815 7.085 0.975 ;
        RECT  6.695 0.430 6.855 2.220 ;
        RECT  6.575 0.770 6.695 1.030 ;
        RECT  3.485 2.060 6.695 2.220 ;
        RECT  6.395 0.310 6.515 0.570 ;
        RECT  6.355 0.310 6.395 0.810 ;
        RECT  6.235 0.410 6.355 0.810 ;
        RECT  6.020 0.650 6.235 0.810 ;
        RECT  0.995 0.310 6.055 0.470 ;
        RECT  5.860 0.650 6.020 1.880 ;
        RECT  4.265 0.650 5.860 0.810 ;
        RECT  4.400 1.720 5.860 1.880 ;
        RECT  3.880 0.675 3.980 0.835 ;
        RECT  3.720 0.675 3.880 1.880 ;
        RECT  3.665 1.605 3.720 1.880 ;
        RECT  3.380 0.650 3.540 1.325 ;
        RECT  3.325 1.565 3.485 2.220 ;
        RECT  1.675 0.650 3.380 0.810 ;
        RECT  3.200 1.565 3.325 1.725 ;
        RECT  3.040 0.990 3.200 1.725 ;
        RECT  2.985 1.905 3.145 2.560 ;
        RECT  2.015 0.990 3.040 1.150 ;
        RECT  2.465 1.905 2.985 2.065 ;
        RECT  2.305 1.905 2.465 2.400 ;
        RECT  1.335 2.240 2.305 2.400 ;
        RECT  1.965 1.675 2.125 1.935 ;
        RECT  1.855 0.990 2.015 1.415 ;
        RECT  1.675 1.675 1.965 1.835 ;
        RECT  1.515 0.650 1.675 1.835 ;
        RECT  1.175 0.695 1.335 2.400 ;
        RECT  0.835 0.310 0.995 1.920 ;
        RECT  0.125 0.715 0.835 0.975 ;
        RECT  0.415 1.760 0.835 1.920 ;
        RECT  0.155 1.760 0.415 2.020 ;
    END
END SDFFHQX4MTH

MACRO SDFFHQX8MTH
    CLASS CORE ;
    FOREIGN SDFFHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.760 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.225 5.890 1.540 ;
        RECT  5.390 1.330 5.495 1.540 ;
        END
        AntennaGateArea 0.1339 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.860 1.030 5.275 1.190 ;
        RECT  4.510 1.030 4.860 1.540 ;
        RECT  4.315 1.030 4.510 1.725 ;
        RECT  4.270 1.465 4.315 1.725 ;
        END
        AntennaGateArea 0.2093 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.865 0.400 14.125 2.380 ;
        RECT  13.105 1.290 13.865 1.665 ;
        RECT  12.845 0.400 13.105 2.380 ;
        END
        AntennaDiffArea 1.164 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.330 3.065 1.620 ;
        END
        AntennaGateArea 0.143 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.305 0.760 1.580 ;
        END
        AntennaGateArea 0.312 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.635 -0.130 14.760 0.130 ;
        RECT  14.375 -0.130 14.635 1.000 ;
        RECT  13.615 -0.130 14.375 0.130 ;
        RECT  13.355 -0.130 13.615 1.000 ;
        RECT  12.595 -0.130 13.355 0.130 ;
        RECT  12.335 -0.130 12.595 1.000 ;
        RECT  11.860 -0.130 12.335 0.130 ;
        RECT  11.260 -0.130 11.860 0.250 ;
        RECT  9.580 -0.130 11.260 0.130 ;
        RECT  9.320 -0.130 9.580 0.250 ;
        RECT  8.695 -0.130 9.320 0.130 ;
        RECT  8.095 -0.130 8.695 0.250 ;
        RECT  0.875 -0.130 8.095 0.130 ;
        RECT  0.615 -0.130 0.875 0.765 ;
        RECT  0.000 -0.130 0.615 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.635 2.740 14.760 3.000 ;
        RECT  14.375 1.785 14.635 3.000 ;
        RECT  13.615 2.740 14.375 3.000 ;
        RECT  13.355 1.885 13.615 3.000 ;
        RECT  12.505 2.740 13.355 3.000 ;
        RECT  11.905 2.415 12.505 3.000 ;
        RECT  9.625 2.740 11.905 3.000 ;
        RECT  9.365 2.620 9.625 3.000 ;
        RECT  8.545 2.740 9.365 3.000 ;
        RECT  8.285 2.620 8.545 3.000 ;
        RECT  3.015 2.740 8.285 3.000 ;
        RECT  2.855 2.245 3.015 3.000 ;
        RECT  2.385 2.740 2.855 3.000 ;
        RECT  2.125 2.620 2.385 3.000 ;
        RECT  0.925 2.740 2.125 3.000 ;
        RECT  0.665 2.105 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.550 1.210 12.600 1.470 ;
        RECT  12.390 1.210 12.550 2.235 ;
        RECT  12.340 1.210 12.390 1.470 ;
        RECT  11.185 2.075 12.390 2.235 ;
        RECT  12.025 1.735 12.135 1.895 ;
        RECT  11.765 0.760 12.025 1.895 ;
        RECT  11.665 1.315 11.765 1.595 ;
        RECT  11.395 1.575 11.445 1.735 ;
        RECT  11.235 0.430 11.395 1.735 ;
        RECT  11.000 0.430 11.235 0.590 ;
        RECT  11.185 1.575 11.235 1.735 ;
        RECT  10.935 1.945 11.185 2.445 ;
        RECT  10.740 0.310 11.000 0.590 ;
        RECT  10.775 0.780 10.935 2.445 ;
        RECT  10.370 0.780 10.775 0.940 ;
        RECT  9.855 2.285 10.775 2.445 ;
        RECT  7.065 0.430 10.740 0.590 ;
        RECT  10.435 1.560 10.595 1.995 ;
        RECT  10.070 1.560 10.435 1.720 ;
        RECT  10.070 0.775 10.120 0.935 ;
        RECT  9.910 0.775 10.070 1.720 ;
        RECT  9.860 0.775 9.910 0.935 ;
        RECT  9.085 1.560 9.910 1.720 ;
        RECT  9.675 1.900 9.855 2.060 ;
        RECT  9.485 1.900 9.675 2.390 ;
        RECT  8.100 2.230 9.485 2.390 ;
        RECT  9.255 1.220 9.290 1.380 ;
        RECT  9.180 1.150 9.255 1.380 ;
        RECT  8.970 0.815 9.180 1.380 ;
        RECT  8.825 1.560 9.085 2.050 ;
        RECT  7.455 0.815 8.970 0.975 ;
        RECT  8.465 1.560 8.825 1.720 ;
        RECT  8.205 1.185 8.465 1.720 ;
        RECT  7.940 2.230 8.100 2.560 ;
        RECT  3.355 2.400 7.940 2.560 ;
        RECT  7.525 1.770 7.785 2.030 ;
        RECT  7.455 1.770 7.525 1.930 ;
        RECT  7.295 0.815 7.455 1.930 ;
        RECT  7.245 0.815 7.295 0.975 ;
        RECT  6.905 0.430 7.065 2.220 ;
        RECT  6.785 0.770 6.905 1.030 ;
        RECT  3.695 2.060 6.905 2.220 ;
        RECT  6.605 0.310 6.725 0.570 ;
        RECT  6.445 0.310 6.605 0.810 ;
        RECT  6.230 0.650 6.445 0.810 ;
        RECT  1.215 0.310 6.265 0.470 ;
        RECT  6.070 0.650 6.230 1.880 ;
        RECT  4.475 0.650 6.070 0.810 ;
        RECT  4.695 1.720 6.070 1.880 ;
        RECT  4.140 0.675 4.190 0.835 ;
        RECT  4.090 0.675 4.140 0.935 ;
        RECT  3.930 0.675 4.090 1.880 ;
        RECT  3.875 1.605 3.930 1.880 ;
        RECT  3.590 0.650 3.750 1.325 ;
        RECT  3.535 1.565 3.695 2.220 ;
        RECT  1.895 0.650 3.590 0.810 ;
        RECT  3.410 1.565 3.535 1.725 ;
        RECT  3.250 0.990 3.410 1.725 ;
        RECT  3.195 1.905 3.355 2.560 ;
        RECT  2.235 0.990 3.250 1.150 ;
        RECT  2.675 1.905 3.195 2.065 ;
        RECT  2.515 1.905 2.675 2.400 ;
        RECT  1.875 2.240 2.515 2.400 ;
        RECT  2.175 1.560 2.335 1.960 ;
        RECT  2.075 0.990 2.235 1.370 ;
        RECT  1.895 1.560 2.175 1.720 ;
        RECT  1.735 0.650 1.895 1.720 ;
        RECT  1.555 1.900 1.875 2.400 ;
        RECT  1.395 0.695 1.555 2.400 ;
        RECT  1.055 0.310 1.215 1.920 ;
        RECT  0.385 0.945 1.055 1.105 ;
        RECT  0.415 1.760 1.055 1.920 ;
        RECT  0.155 1.760 0.415 2.020 ;
        RECT  0.125 0.705 0.385 1.105 ;
    END
END SDFFHQX8MTH

MACRO SDFFHX1MTH
    CLASS CORE ;
    FOREIGN SDFFHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.120 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.450 0.990 5.610 1.350 ;
        RECT  4.450 0.990 5.450 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.1131 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.810 0.765 13.020 1.995 ;
        RECT  12.735 0.765 12.810 1.025 ;
        RECT  12.705 1.735 12.810 1.995 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.580 0.815 11.790 1.995 ;
        END
        AntennaDiffArea 0.29 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.330 2.575 1.620 ;
        END
        AntennaGateArea 0.0663 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.355 1.990 ;
        END
        AntennaGateArea 0.1365 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.795 -0.130 13.120 0.130 ;
        RECT  12.515 -0.130 12.795 0.300 ;
        RECT  12.320 -0.130 12.515 0.130 ;
        RECT  11.820 -0.130 12.320 0.300 ;
        RECT  10.900 -0.130 11.820 0.130 ;
        RECT  10.740 -0.130 10.900 0.620 ;
        RECT  9.150 -0.130 10.740 0.130 ;
        RECT  8.890 -0.130 9.150 0.250 ;
        RECT  7.990 -0.130 8.890 0.130 ;
        RECT  7.730 -0.130 7.990 0.250 ;
        RECT  0.355 -0.130 7.730 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.670 2.740 13.120 3.000 ;
        RECT  12.170 2.570 12.670 3.000 ;
        RECT  11.060 2.740 12.170 3.000 ;
        RECT  10.900 2.230 11.060 3.000 ;
        RECT  8.640 2.740 10.900 3.000 ;
        RECT  8.040 2.205 8.640 3.000 ;
        RECT  7.075 2.740 8.040 3.000 ;
        RECT  6.815 2.570 7.075 3.000 ;
        RECT  2.695 2.740 6.815 3.000 ;
        RECT  2.535 2.150 2.695 3.000 ;
        RECT  0.905 2.740 2.535 3.000 ;
        RECT  0.745 2.570 0.905 3.000 ;
        RECT  0.000 2.740 0.745 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.130 1.250 12.575 1.510 ;
        RECT  11.970 1.250 12.130 2.335 ;
        RECT  11.810 2.175 11.970 2.335 ;
        RECT  11.550 2.175 11.810 2.560 ;
        RECT  11.400 2.175 11.550 2.335 ;
        RECT  11.400 0.355 11.520 0.565 ;
        RECT  11.240 0.355 11.400 2.335 ;
        RECT  10.870 1.265 11.240 1.525 ;
        RECT  10.350 2.400 10.720 2.560 ;
        RECT  10.540 0.810 10.600 1.710 ;
        RECT  10.440 0.430 10.540 1.710 ;
        RECT  10.380 0.430 10.440 0.975 ;
        RECT  10.030 0.430 10.380 0.590 ;
        RECT  10.250 1.940 10.350 2.560 ;
        RECT  10.200 1.185 10.250 2.560 ;
        RECT  10.090 0.815 10.200 2.560 ;
        RECT  10.040 0.815 10.090 1.345 ;
        RECT  9.940 0.815 10.040 0.975 ;
        RECT  9.770 0.345 10.030 0.590 ;
        RECT  9.720 1.840 9.790 2.100 ;
        RECT  8.550 0.430 9.770 0.590 ;
        RECT  9.560 0.800 9.720 2.100 ;
        RECT  9.110 2.385 9.580 2.545 ;
        RECT  9.430 0.800 9.560 0.960 ;
        RECT  9.290 1.525 9.560 2.100 ;
        RECT  9.180 1.185 9.350 1.345 ;
        RECT  8.090 1.525 9.290 1.685 ;
        RECT  9.020 0.820 9.180 1.345 ;
        RECT  8.950 1.865 9.110 2.545 ;
        RECT  8.350 0.820 9.020 0.980 ;
        RECT  7.780 1.865 8.950 2.025 ;
        RECT  8.290 0.310 8.550 0.590 ;
        RECT  8.090 0.770 8.350 0.980 ;
        RECT  7.425 0.430 8.290 0.590 ;
        RECT  7.080 0.820 8.090 0.980 ;
        RECT  7.930 1.195 8.090 1.685 ;
        RECT  7.830 1.195 7.930 1.355 ;
        RECT  7.620 1.865 7.780 2.560 ;
        RECT  7.520 2.130 7.620 2.560 ;
        RECT  6.635 2.130 7.520 2.290 ;
        RECT  7.265 0.380 7.425 0.590 ;
        RECT  7.080 1.690 7.355 1.950 ;
        RECT  6.740 0.380 7.265 0.540 ;
        RECT  6.920 0.720 7.080 1.950 ;
        RECT  6.580 0.380 6.740 1.550 ;
        RECT  6.475 2.130 6.635 2.560 ;
        RECT  6.325 0.750 6.580 1.550 ;
        RECT  3.035 2.400 6.475 2.560 ;
        RECT  6.240 0.310 6.400 0.570 ;
        RECT  6.295 1.290 6.325 1.550 ;
        RECT  6.135 1.290 6.295 2.220 ;
        RECT  6.145 0.410 6.240 0.570 ;
        RECT  5.985 0.410 6.145 0.810 ;
        RECT  3.375 2.060 6.135 2.220 ;
        RECT  5.950 0.650 5.985 0.810 ;
        RECT  5.790 0.650 5.950 1.880 ;
        RECT  0.695 0.310 5.805 0.470 ;
        RECT  4.005 0.650 5.790 0.810 ;
        RECT  4.125 1.720 5.790 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.435 0.650 3.555 0.810 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.095 0.650 3.255 1.230 ;
        RECT  2.915 1.465 3.215 1.625 ;
        RECT  1.035 0.650 3.095 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.755 0.990 2.915 1.625 ;
        RECT  1.615 1.805 2.875 1.965 ;
        RECT  1.735 0.990 2.755 1.150 ;
        RECT  1.965 2.145 2.125 2.510 ;
        RECT  1.275 2.350 1.965 2.510 ;
        RECT  1.575 0.990 1.735 1.625 ;
        RECT  1.455 1.805 1.615 2.170 ;
        RECT  1.375 1.805 1.455 1.965 ;
        RECT  1.215 0.990 1.375 1.965 ;
        RECT  1.115 2.145 1.275 2.510 ;
        RECT  1.035 2.145 1.115 2.305 ;
        RECT  0.875 0.650 1.035 2.305 ;
        RECT  0.535 0.310 0.695 2.345 ;
        RECT  0.125 0.765 0.535 1.025 ;
        RECT  0.385 2.185 0.535 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFHX1MTH

MACRO SDFFHX2MTH
    CLASS CORE ;
    FOREIGN SDFFHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.450 0.990 5.610 1.350 ;
        RECT  4.450 0.990 5.450 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.1274 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.175 0.765 13.430 1.950 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.160 1.290 12.200 1.580 ;
        RECT  12.050 0.425 12.160 1.580 ;
        RECT  11.890 0.425 12.050 1.985 ;
        END
        AntennaDiffArea 0.417 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.330 2.575 1.620 ;
        END
        AntennaGateArea 0.0923 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.355 1.910 ;
        END
        AntennaGateArea 0.1456 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.040 -0.130 13.530 0.130 ;
        RECT  12.700 -0.130 13.040 0.300 ;
        RECT  12.440 -0.130 12.700 1.025 ;
        RECT  10.950 -0.130 12.440 0.130 ;
        RECT  10.690 -0.130 10.950 0.250 ;
        RECT  9.150 -0.130 10.690 0.130 ;
        RECT  8.890 -0.130 9.150 0.250 ;
        RECT  7.990 -0.130 8.890 0.130 ;
        RECT  7.730 -0.130 7.990 0.250 ;
        RECT  0.355 -0.130 7.730 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.040 2.740 13.530 3.000 ;
        RECT  12.780 2.190 13.040 3.000 ;
        RECT  12.440 2.570 12.780 3.000 ;
        RECT  11.350 2.740 12.440 3.000 ;
        RECT  11.190 2.235 11.350 3.000 ;
        RECT  8.150 2.740 11.190 3.000 ;
        RECT  7.890 2.620 8.150 3.000 ;
        RECT  2.695 2.740 7.890 3.000 ;
        RECT  2.535 2.150 2.695 3.000 ;
        RECT  0.690 2.740 2.535 3.000 ;
        RECT  0.430 2.570 0.690 3.000 ;
        RECT  0.000 2.740 0.430 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.705 1.250 12.965 1.510 ;
        RECT  12.540 1.350 12.705 1.510 ;
        RECT  12.380 1.350 12.540 2.325 ;
        RECT  12.130 2.165 12.380 2.325 ;
        RECT  11.870 2.165 12.130 2.515 ;
        RECT  11.690 2.165 11.870 2.325 ;
        RECT  11.530 1.265 11.690 2.325 ;
        RECT  11.520 1.265 11.530 1.525 ;
        RECT  11.260 0.440 11.520 1.525 ;
        RECT  11.190 1.265 11.260 1.525 ;
        RECT  10.710 2.400 11.010 2.560 ;
        RECT  10.760 0.435 10.920 1.710 ;
        RECT  10.460 0.435 10.760 0.595 ;
        RECT  10.500 1.940 10.710 2.560 ;
        RECT  10.490 1.940 10.500 2.100 ;
        RECT  9.810 2.400 10.500 2.560 ;
        RECT  10.330 0.815 10.490 2.100 ;
        RECT  10.200 0.310 10.460 0.595 ;
        RECT  9.940 0.815 10.330 0.975 ;
        RECT  8.550 0.435 10.200 0.595 ;
        RECT  9.990 1.525 10.150 2.075 ;
        RECT  9.720 1.525 9.990 1.685 ;
        RECT  9.650 1.865 9.810 2.560 ;
        RECT  9.560 0.800 9.720 1.685 ;
        RECT  9.350 1.865 9.650 2.025 ;
        RECT  9.430 0.800 9.560 0.960 ;
        RECT  8.700 1.525 9.560 1.685 ;
        RECT  9.210 2.230 9.470 2.545 ;
        RECT  9.180 1.185 9.350 1.345 ;
        RECT  7.710 2.230 9.210 2.390 ;
        RECT  9.020 0.820 9.180 1.345 ;
        RECT  7.080 0.820 9.020 0.980 ;
        RECT  8.440 1.525 8.700 2.050 ;
        RECT  8.290 0.325 8.550 0.595 ;
        RECT  8.090 1.525 8.440 1.685 ;
        RECT  7.425 0.435 8.290 0.595 ;
        RECT  7.930 1.195 8.090 1.685 ;
        RECT  7.830 1.195 7.930 1.355 ;
        RECT  7.450 2.230 7.710 2.560 ;
        RECT  3.035 2.400 7.450 2.560 ;
        RECT  7.265 0.380 7.425 0.595 ;
        RECT  6.740 0.380 7.265 0.540 ;
        RECT  7.080 1.690 7.255 1.950 ;
        RECT  6.920 0.720 7.080 1.950 ;
        RECT  6.580 0.380 6.740 0.910 ;
        RECT  6.555 0.750 6.580 0.910 ;
        RECT  6.395 0.750 6.555 2.220 ;
        RECT  6.240 0.310 6.400 0.570 ;
        RECT  6.325 0.750 6.395 1.010 ;
        RECT  3.375 2.060 6.395 2.220 ;
        RECT  6.145 0.410 6.240 0.570 ;
        RECT  5.985 0.410 6.145 0.810 ;
        RECT  5.950 0.650 5.985 0.810 ;
        RECT  5.790 0.650 5.950 1.880 ;
        RECT  0.695 0.310 5.805 0.470 ;
        RECT  4.005 0.650 5.790 0.810 ;
        RECT  4.125 1.720 5.790 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.435 0.650 3.555 0.810 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.095 0.650 3.255 1.230 ;
        RECT  2.915 1.465 3.215 1.625 ;
        RECT  1.035 0.650 3.095 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.755 0.990 2.915 1.625 ;
        RECT  1.665 1.805 2.875 1.965 ;
        RECT  1.735 0.990 2.755 1.150 ;
        RECT  1.965 2.145 2.125 2.465 ;
        RECT  1.035 2.305 1.965 2.465 ;
        RECT  1.575 0.990 1.735 1.625 ;
        RECT  1.405 1.805 1.665 2.120 ;
        RECT  1.375 1.805 1.405 1.965 ;
        RECT  1.215 0.990 1.375 1.965 ;
        RECT  0.875 0.650 1.035 2.465 ;
        RECT  0.535 0.310 0.695 2.250 ;
        RECT  0.125 0.765 0.535 1.025 ;
        RECT  0.385 2.090 0.535 2.250 ;
        RECT  0.125 2.090 0.385 2.325 ;
    END
END SDFFHX2MTH

MACRO SDFFHX4MTH
    CLASS CORE ;
    FOREIGN SDFFHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.940 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.0832 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 0.990 5.515 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.182 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.630 0.765 13.840 1.945 ;
        RECT  13.555 0.765 13.630 1.025 ;
        RECT  13.555 1.685 13.630 1.945 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.835 1.290 13.020 1.580 ;
        RECT  12.580 0.425 12.835 1.945 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.330 2.575 1.620 ;
        END
        AntennaGateArea 0.1586 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.355 1.990 ;
        END
        AntennaGateArea 0.2041 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.375 -0.130 13.940 0.130 ;
        RECT  13.115 -0.130 13.375 0.570 ;
        RECT  12.325 -0.130 13.115 0.130 ;
        RECT  12.065 -0.130 12.325 1.020 ;
        RECT  11.195 -0.130 12.065 0.130 ;
        RECT  11.035 -0.130 11.195 0.730 ;
        RECT  9.175 -0.130 11.035 0.130 ;
        RECT  8.915 -0.130 9.175 0.250 ;
        RECT  8.015 -0.130 8.915 0.130 ;
        RECT  7.755 -0.130 8.015 0.250 ;
        RECT  0.355 -0.130 7.755 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.375 2.740 13.940 3.000 ;
        RECT  13.115 2.465 13.375 3.000 ;
        RECT  12.295 2.740 13.115 3.000 ;
        RECT  12.035 2.465 12.295 3.000 ;
        RECT  11.675 2.740 12.035 3.000 ;
        RECT  11.415 2.465 11.675 3.000 ;
        RECT  8.175 2.740 11.415 3.000 ;
        RECT  7.915 2.620 8.175 3.000 ;
        RECT  2.695 2.740 7.915 3.000 ;
        RECT  2.535 2.150 2.695 3.000 ;
        RECT  0.000 2.740 2.535 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.370 1.245 13.450 1.505 ;
        RECT  13.210 1.245 13.370 2.285 ;
        RECT  12.385 2.125 13.210 2.285 ;
        RECT  12.225 1.785 12.385 2.285 ;
        RECT  11.845 1.785 12.225 1.945 ;
        RECT  10.735 2.125 12.045 2.285 ;
        RECT  11.815 1.685 11.845 1.945 ;
        RECT  11.585 0.490 11.815 1.945 ;
        RECT  11.555 0.490 11.585 1.400 ;
        RECT  11.215 1.135 11.555 1.400 ;
        RECT  10.855 1.450 10.945 1.710 ;
        RECT  10.695 0.430 10.855 1.710 ;
        RECT  10.515 1.900 10.735 2.560 ;
        RECT  10.485 0.430 10.695 0.590 ;
        RECT  10.355 0.815 10.515 2.560 ;
        RECT  10.225 0.310 10.485 0.590 ;
        RECT  9.965 0.815 10.355 0.975 ;
        RECT  9.835 2.400 10.355 2.560 ;
        RECT  8.575 0.430 10.225 0.590 ;
        RECT  10.015 1.525 10.175 2.075 ;
        RECT  9.745 1.525 10.015 1.720 ;
        RECT  9.675 1.900 9.835 2.560 ;
        RECT  9.585 0.800 9.745 1.720 ;
        RECT  9.375 1.900 9.675 2.060 ;
        RECT  9.455 0.800 9.585 0.960 ;
        RECT  8.725 1.560 9.585 1.720 ;
        RECT  9.235 2.280 9.495 2.545 ;
        RECT  9.205 1.220 9.375 1.380 ;
        RECT  7.735 2.280 9.235 2.440 ;
        RECT  9.115 0.815 9.205 1.380 ;
        RECT  9.045 0.815 9.115 1.370 ;
        RECT  7.335 0.815 9.045 0.975 ;
        RECT  8.465 1.560 8.725 2.050 ;
        RECT  8.315 0.325 8.575 0.590 ;
        RECT  8.115 1.560 8.465 1.720 ;
        RECT  7.450 0.430 8.315 0.590 ;
        RECT  7.955 1.195 8.115 1.720 ;
        RECT  7.855 1.195 7.955 1.355 ;
        RECT  7.475 2.280 7.735 2.560 ;
        RECT  3.035 2.400 7.475 2.560 ;
        RECT  7.290 0.310 7.450 0.590 ;
        RECT  7.175 0.815 7.335 1.950 ;
        RECT  6.765 0.310 7.290 0.470 ;
        RECT  7.105 0.815 7.175 0.980 ;
        RECT  6.945 0.720 7.105 0.980 ;
        RECT  6.685 0.310 6.765 0.910 ;
        RECT  6.605 0.310 6.685 2.220 ;
        RECT  6.525 0.750 6.605 2.220 ;
        RECT  6.325 0.750 6.525 1.010 ;
        RECT  3.375 2.060 6.525 2.220 ;
        RECT  6.145 0.310 6.425 0.470 ;
        RECT  5.985 0.310 6.145 0.810 ;
        RECT  5.950 0.650 5.985 0.810 ;
        RECT  5.790 0.650 5.950 1.880 ;
        RECT  0.695 0.310 5.805 0.470 ;
        RECT  3.945 0.650 5.790 0.810 ;
        RECT  4.095 1.720 5.790 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.435 0.650 3.555 0.810 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.095 0.650 3.255 1.230 ;
        RECT  2.915 1.465 3.215 1.625 ;
        RECT  1.035 0.650 3.095 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.755 0.990 2.915 1.625 ;
        RECT  1.665 1.805 2.875 1.965 ;
        RECT  1.735 0.990 2.755 1.150 ;
        RECT  1.965 2.145 2.125 2.465 ;
        RECT  1.035 2.305 1.965 2.465 ;
        RECT  1.575 0.990 1.735 1.625 ;
        RECT  1.405 1.805 1.665 2.120 ;
        RECT  1.375 1.805 1.405 1.965 ;
        RECT  1.215 0.990 1.375 1.965 ;
        RECT  0.875 0.650 1.035 2.465 ;
        RECT  0.535 0.310 0.695 2.345 ;
        RECT  0.125 0.765 0.535 1.025 ;
        RECT  0.385 2.185 0.535 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFHX4MTH

MACRO SDFFHX8MTH
    CLASS CORE ;
    FOREIGN SDFFHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.760 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.0832 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 0.990 5.515 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.182 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.450 0.765 14.660 1.945 ;
        RECT  14.375 0.765 14.450 1.025 ;
        RECT  14.375 1.685 14.450 1.945 ;
        END
        AntennaDiffArea 0.209 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.410 0.425 13.665 1.945 ;
        RECT  12.735 1.290 13.410 1.580 ;
        RECT  12.480 0.425 12.735 1.945 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 1.330 2.575 1.620 ;
        END
        AntennaGateArea 0.1586 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.355 1.990 ;
        END
        AntennaGateArea 0.2041 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.205 -0.130 14.760 0.130 ;
        RECT  13.945 -0.130 14.205 0.570 ;
        RECT  12.195 -0.130 13.945 0.130 ;
        RECT  11.935 -0.130 12.195 0.385 ;
        RECT  11.195 -0.130 11.935 0.130 ;
        RECT  11.035 -0.130 11.195 0.730 ;
        RECT  9.175 -0.130 11.035 0.130 ;
        RECT  8.915 -0.130 9.175 0.250 ;
        RECT  8.015 -0.130 8.915 0.130 ;
        RECT  7.755 -0.130 8.015 0.250 ;
        RECT  0.355 -0.130 7.755 0.130 ;
        RECT  0.195 -0.130 0.355 0.300 ;
        RECT  0.000 -0.130 0.195 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.205 2.740 14.760 3.000 ;
        RECT  13.945 2.465 14.205 3.000 ;
        RECT  12.125 2.740 13.945 3.000 ;
        RECT  11.525 2.530 12.125 3.000 ;
        RECT  8.175 2.740 11.525 3.000 ;
        RECT  7.915 2.620 8.175 3.000 ;
        RECT  2.695 2.740 7.915 3.000 ;
        RECT  2.535 2.150 2.695 3.000 ;
        RECT  0.000 2.740 2.535 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.190 1.245 14.270 1.505 ;
        RECT  14.030 1.245 14.190 2.285 ;
        RECT  12.285 2.125 14.030 2.285 ;
        RECT  12.125 1.785 12.285 2.285 ;
        RECT  11.815 1.785 12.125 1.945 ;
        RECT  10.735 2.125 11.945 2.285 ;
        RECT  11.555 0.685 11.815 1.945 ;
        RECT  11.485 1.310 11.555 1.945 ;
        RECT  11.215 1.310 11.485 1.575 ;
        RECT  10.855 1.625 10.945 1.885 ;
        RECT  10.695 0.430 10.855 1.885 ;
        RECT  10.515 2.125 10.735 2.560 ;
        RECT  10.485 0.430 10.695 0.590 ;
        RECT  10.355 0.815 10.515 2.560 ;
        RECT  10.225 0.310 10.485 0.590 ;
        RECT  9.965 0.815 10.355 0.975 ;
        RECT  9.835 2.400 10.355 2.560 ;
        RECT  8.575 0.430 10.225 0.590 ;
        RECT  10.015 1.525 10.175 2.075 ;
        RECT  9.745 1.525 10.015 1.720 ;
        RECT  9.675 1.900 9.835 2.560 ;
        RECT  9.585 0.800 9.745 1.720 ;
        RECT  9.375 1.900 9.675 2.060 ;
        RECT  9.455 0.800 9.585 0.960 ;
        RECT  8.725 1.560 9.585 1.720 ;
        RECT  9.235 2.280 9.495 2.545 ;
        RECT  9.205 1.220 9.375 1.380 ;
        RECT  7.735 2.280 9.235 2.440 ;
        RECT  9.115 0.815 9.205 1.380 ;
        RECT  9.045 0.815 9.115 1.370 ;
        RECT  7.335 0.815 9.045 0.975 ;
        RECT  8.465 1.560 8.725 2.050 ;
        RECT  8.315 0.325 8.575 0.590 ;
        RECT  8.115 1.560 8.465 1.720 ;
        RECT  7.450 0.430 8.315 0.590 ;
        RECT  7.955 1.195 8.115 1.720 ;
        RECT  7.855 1.195 7.955 1.355 ;
        RECT  7.475 2.280 7.735 2.560 ;
        RECT  3.035 2.400 7.475 2.560 ;
        RECT  7.290 0.310 7.450 0.590 ;
        RECT  7.175 0.815 7.335 1.950 ;
        RECT  6.765 0.310 7.290 0.470 ;
        RECT  7.105 0.815 7.175 0.980 ;
        RECT  6.945 0.720 7.105 0.980 ;
        RECT  6.685 0.310 6.765 0.910 ;
        RECT  6.605 0.310 6.685 2.220 ;
        RECT  6.525 0.750 6.605 2.220 ;
        RECT  6.325 0.750 6.525 1.010 ;
        RECT  3.375 2.060 6.525 2.220 ;
        RECT  6.145 0.310 6.425 0.470 ;
        RECT  5.985 0.310 6.145 0.810 ;
        RECT  5.950 0.650 5.985 0.810 ;
        RECT  5.790 0.650 5.950 1.880 ;
        RECT  0.695 0.310 5.805 0.470 ;
        RECT  3.945 0.650 5.790 0.810 ;
        RECT  4.095 1.720 5.790 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.435 0.650 3.555 0.810 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.095 0.650 3.255 1.230 ;
        RECT  2.915 1.465 3.215 1.625 ;
        RECT  1.035 0.650 3.095 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.755 0.990 2.915 1.625 ;
        RECT  1.665 1.805 2.875 1.965 ;
        RECT  1.735 0.990 2.755 1.150 ;
        RECT  1.965 2.145 2.125 2.465 ;
        RECT  1.035 2.305 1.965 2.465 ;
        RECT  1.575 0.990 1.735 1.625 ;
        RECT  1.405 1.805 1.665 2.120 ;
        RECT  1.375 1.805 1.405 1.965 ;
        RECT  1.215 0.990 1.375 1.965 ;
        RECT  0.875 0.650 1.035 2.465 ;
        RECT  0.535 0.310 0.695 2.345 ;
        RECT  0.125 0.765 0.535 1.025 ;
        RECT  0.385 2.185 0.535 2.345 ;
        RECT  0.125 2.185 0.385 2.445 ;
    END
END SDFFHX8MTH

MACRO SDFFNHX1MTH
    CLASS CORE ;
    FOREIGN SDFFNHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.440 0.990 5.600 1.260 ;
        RECT  4.450 0.990 5.440 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.270 0.765 13.430 1.990 ;
        RECT  13.145 0.765 13.270 1.025 ;
        RECT  13.145 1.700 13.270 1.990 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.415 1.290 12.610 1.580 ;
        RECT  12.255 0.730 12.415 1.955 ;
        RECT  12.125 0.730 12.255 0.990 ;
        END
        AntennaDiffArea 0.274 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.580 1.590 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.240 0.430 1.710 ;
        END
        AntennaGateArea 0.1378 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.095 -0.130 13.530 0.130 ;
        RECT  12.155 -0.130 13.095 0.340 ;
        RECT  11.205 -0.130 12.155 0.130 ;
        RECT  10.605 -0.130 11.205 0.300 ;
        RECT  9.475 -0.130 10.605 0.130 ;
        RECT  8.875 -0.130 9.475 0.250 ;
        RECT  8.255 -0.130 8.875 0.130 ;
        RECT  7.655 -0.130 8.255 0.250 ;
        RECT  0.430 -0.130 7.655 0.130 ;
        RECT  0.270 -0.130 0.430 0.350 ;
        RECT  0.000 -0.130 0.270 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.005 2.740 13.530 3.000 ;
        RECT  12.745 2.505 13.005 3.000 ;
        RECT  11.735 2.740 12.745 3.000 ;
        RECT  11.575 1.795 11.735 3.000 ;
        RECT  9.235 2.740 11.575 3.000 ;
        RECT  8.635 2.620 9.235 3.000 ;
        RECT  6.935 2.740 8.635 3.000 ;
        RECT  6.675 2.560 6.935 3.000 ;
        RECT  2.695 2.740 6.675 3.000 ;
        RECT  2.535 2.145 2.695 3.000 ;
        RECT  0.770 2.740 2.535 3.000 ;
        RECT  0.170 2.505 0.770 3.000 ;
        RECT  0.000 2.740 0.170 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.955 1.250 13.080 1.510 ;
        RECT  12.795 1.250 12.955 2.325 ;
        RECT  12.385 2.165 12.795 2.325 ;
        RECT  12.125 2.165 12.385 2.430 ;
        RECT  12.075 2.165 12.125 2.325 ;
        RECT  11.915 1.365 12.075 2.325 ;
        RECT  11.775 1.365 11.915 1.580 ;
        RECT  11.775 0.550 11.875 0.710 ;
        RECT  11.615 0.550 11.775 1.580 ;
        RECT  11.315 1.320 11.615 1.580 ;
        RECT  10.885 0.480 11.050 1.750 ;
        RECT  10.140 0.480 10.885 0.640 ;
        RECT  10.700 2.400 10.800 2.560 ;
        RECT  10.540 0.820 10.700 2.560 ;
        RECT  10.050 0.820 10.540 0.980 ;
        RECT  10.195 1.400 10.355 2.475 ;
        RECT  9.575 2.315 10.195 2.475 ;
        RECT  9.880 0.380 10.140 0.640 ;
        RECT  9.870 1.960 10.015 2.135 ;
        RECT  8.695 0.480 9.880 0.640 ;
        RECT  9.755 0.820 9.870 2.135 ;
        RECT  9.710 0.820 9.755 2.100 ;
        RECT  9.540 0.820 9.710 0.980 ;
        RECT  8.880 1.940 9.710 2.100 ;
        RECT  9.415 2.280 9.575 2.475 ;
        RECT  9.270 1.590 9.530 1.750 ;
        RECT  8.400 2.280 9.415 2.440 ;
        RECT  9.110 0.820 9.270 1.750 ;
        RECT  8.200 0.820 9.110 0.980 ;
        RECT  8.620 1.280 8.880 2.100 ;
        RECT  8.485 0.405 8.695 0.640 ;
        RECT  8.435 0.405 8.485 0.595 ;
        RECT  6.885 0.435 8.435 0.595 ;
        RECT  8.140 2.280 8.400 2.485 ;
        RECT  8.040 0.775 8.200 2.085 ;
        RECT  7.420 2.280 8.140 2.440 ;
        RECT  7.225 0.775 8.040 0.935 ;
        RECT  7.600 1.925 8.040 2.085 ;
        RECT  7.260 1.215 7.420 2.440 ;
        RECT  6.765 1.215 7.260 1.375 ;
        RECT  6.355 2.220 7.260 2.380 ;
        RECT  7.065 0.775 7.225 1.035 ;
        RECT  6.325 1.555 7.080 1.715 ;
        RECT  6.725 0.435 6.885 0.810 ;
        RECT  6.505 0.990 6.765 1.375 ;
        RECT  6.325 0.650 6.725 0.810 ;
        RECT  5.985 0.310 6.545 0.470 ;
        RECT  6.195 2.220 6.355 2.560 ;
        RECT  6.165 0.650 6.325 1.940 ;
        RECT  3.035 2.400 6.195 2.560 ;
        RECT  5.950 1.780 6.165 1.940 ;
        RECT  5.825 0.310 5.985 1.600 ;
        RECT  5.790 1.780 5.950 2.220 ;
        RECT  4.120 0.650 5.825 0.810 ;
        RECT  5.610 1.440 5.825 1.600 ;
        RECT  3.375 2.060 5.790 2.220 ;
        RECT  0.770 0.310 5.645 0.470 ;
        RECT  5.450 1.440 5.610 1.880 ;
        RECT  4.125 1.720 5.450 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.440 0.650 3.555 0.810 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.260 0.970 3.355 1.230 ;
        RECT  3.100 0.650 3.260 1.230 ;
        RECT  2.920 1.465 3.215 1.625 ;
        RECT  1.110 0.650 3.100 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.760 0.990 2.920 1.625 ;
        RECT  1.980 1.805 2.875 1.965 ;
        RECT  1.450 0.990 2.760 1.150 ;
        RECT  1.965 2.145 2.125 2.560 ;
        RECT  1.820 1.720 1.980 1.965 ;
        RECT  1.110 2.400 1.965 2.560 ;
        RECT  1.790 1.720 1.820 1.880 ;
        RECT  1.630 1.620 1.790 1.880 ;
        RECT  1.450 2.060 1.665 2.220 ;
        RECT  1.290 0.990 1.450 2.220 ;
        RECT  0.950 0.650 1.110 2.560 ;
        RECT  0.610 0.310 0.770 2.170 ;
        RECT  0.125 0.765 0.610 1.025 ;
        RECT  0.385 1.980 0.610 2.170 ;
        RECT  0.125 1.980 0.385 2.240 ;
    END
END SDFFNHX1MTH

MACRO SDFFNHX2MTH
    CLASS CORE ;
    FOREIGN SDFFNHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.940 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.450 0.990 5.610 1.260 ;
        RECT  4.450 0.990 5.450 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.680 0.765 13.840 1.990 ;
        RECT  13.555 0.765 13.680 1.025 ;
        RECT  13.555 1.700 13.680 1.990 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.825 1.290 13.020 1.580 ;
        RECT  12.665 0.380 12.825 1.985 ;
        RECT  12.535 0.380 12.665 0.980 ;
        END
        AntennaDiffArea 0.437 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.580 1.590 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.240 0.430 1.710 ;
        END
        AntennaGateArea 0.1378 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.675 -0.130 13.940 0.130 ;
        RECT  13.075 -0.130 13.675 0.515 ;
        RECT  11.840 -0.130 13.075 0.130 ;
        RECT  11.240 -0.130 11.840 0.300 ;
        RECT  9.650 -0.130 11.240 0.130 ;
        RECT  9.390 -0.130 9.650 0.300 ;
        RECT  8.480 -0.130 9.390 0.130 ;
        RECT  8.220 -0.130 8.480 0.250 ;
        RECT  0.430 -0.130 8.220 0.130 ;
        RECT  0.270 -0.130 0.430 0.330 ;
        RECT  0.000 -0.130 0.270 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.755 2.740 13.940 3.000 ;
        RECT  13.155 2.515 13.755 3.000 ;
        RECT  12.145 2.740 13.155 3.000 ;
        RECT  11.985 1.795 12.145 3.000 ;
        RECT  9.885 2.740 11.985 3.000 ;
        RECT  9.285 2.595 9.885 3.000 ;
        RECT  7.290 2.740 9.285 3.000 ;
        RECT  7.030 2.280 7.290 3.000 ;
        RECT  2.695 2.740 7.030 3.000 ;
        RECT  2.535 2.145 2.695 3.000 ;
        RECT  0.765 2.740 2.535 3.000 ;
        RECT  0.605 2.505 0.765 3.000 ;
        RECT  0.000 2.740 0.605 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.365 1.250 13.490 1.510 ;
        RECT  13.205 1.250 13.365 2.325 ;
        RECT  12.795 2.165 13.205 2.325 ;
        RECT  12.535 2.165 12.795 2.520 ;
        RECT  12.485 2.165 12.535 2.325 ;
        RECT  12.325 1.415 12.485 2.325 ;
        RECT  12.185 1.415 12.325 1.580 ;
        RECT  12.185 0.550 12.285 0.710 ;
        RECT  12.025 0.550 12.185 1.580 ;
        RECT  11.725 1.320 12.025 1.580 ;
        RECT  11.295 0.480 11.455 1.750 ;
        RECT  10.960 0.480 11.295 0.640 ;
        RECT  11.110 2.400 11.210 2.560 ;
        RECT  10.950 0.820 11.110 2.560 ;
        RECT  10.700 0.310 10.960 0.640 ;
        RECT  10.440 0.820 10.950 0.980 ;
        RECT  10.605 1.375 10.765 2.410 ;
        RECT  9.050 0.480 10.700 0.640 ;
        RECT  8.950 2.250 10.605 2.410 ;
        RECT  10.190 1.910 10.425 2.070 ;
        RECT  10.030 0.820 10.190 2.070 ;
        RECT  9.930 0.820 10.030 0.980 ;
        RECT  9.290 1.910 10.030 2.070 ;
        RECT  9.680 1.295 9.850 1.555 ;
        RECT  9.520 0.850 9.680 1.555 ;
        RECT  8.610 0.850 9.520 1.010 ;
        RECT  9.030 1.490 9.290 2.070 ;
        RECT  8.790 0.435 9.050 0.640 ;
        RECT  8.790 2.250 8.950 2.440 ;
        RECT  7.240 0.435 8.790 0.595 ;
        RECT  7.830 2.280 8.790 2.440 ;
        RECT  8.450 0.775 8.610 2.070 ;
        RECT  7.580 0.775 8.450 0.935 ;
        RECT  8.010 1.910 8.450 2.070 ;
        RECT  7.670 1.215 7.830 2.440 ;
        RECT  6.990 1.215 7.670 1.375 ;
        RECT  6.850 1.940 7.670 2.100 ;
        RECT  7.420 0.775 7.580 1.035 ;
        RECT  6.550 1.555 7.490 1.715 ;
        RECT  7.080 0.435 7.240 0.810 ;
        RECT  6.550 0.650 7.080 0.810 ;
        RECT  6.730 0.990 6.990 1.375 ;
        RECT  6.210 0.310 6.900 0.470 ;
        RECT  6.690 1.940 6.850 2.280 ;
        RECT  6.290 2.120 6.690 2.280 ;
        RECT  6.510 0.650 6.550 1.715 ;
        RECT  6.390 0.650 6.510 1.940 ;
        RECT  6.350 1.555 6.390 1.940 ;
        RECT  5.950 1.780 6.350 1.940 ;
        RECT  6.130 2.120 6.290 2.560 ;
        RECT  6.170 0.310 6.210 0.810 ;
        RECT  6.050 0.310 6.170 1.600 ;
        RECT  3.035 2.400 6.130 2.560 ;
        RECT  6.010 0.650 6.050 1.600 ;
        RECT  4.120 0.650 6.010 0.810 ;
        RECT  5.610 1.440 6.010 1.600 ;
        RECT  5.790 1.780 5.950 2.220 ;
        RECT  0.770 0.310 5.870 0.470 ;
        RECT  3.375 2.060 5.790 2.220 ;
        RECT  5.450 1.440 5.610 1.880 ;
        RECT  4.125 1.720 5.450 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.440 0.650 3.555 0.810 ;
        RECT  3.260 0.990 3.375 1.250 ;
        RECT  3.215 1.465 3.375 2.220 ;
        RECT  3.100 0.650 3.260 1.250 ;
        RECT  2.920 1.465 3.215 1.625 ;
        RECT  1.110 0.650 3.100 0.810 ;
        RECT  2.875 1.805 3.035 2.560 ;
        RECT  2.760 0.990 2.920 1.625 ;
        RECT  1.980 1.805 2.875 1.965 ;
        RECT  1.450 0.990 2.760 1.150 ;
        RECT  1.965 2.145 2.125 2.560 ;
        RECT  1.820 1.720 1.980 1.965 ;
        RECT  1.110 2.400 1.965 2.560 ;
        RECT  1.790 1.720 1.820 1.880 ;
        RECT  1.630 1.620 1.790 1.880 ;
        RECT  1.450 2.060 1.665 2.220 ;
        RECT  1.290 0.990 1.450 2.220 ;
        RECT  0.950 0.650 1.110 2.560 ;
        RECT  0.610 0.310 0.770 2.170 ;
        RECT  0.125 0.765 0.610 1.025 ;
        RECT  0.385 2.010 0.610 2.170 ;
        RECT  0.125 2.010 0.385 2.270 ;
    END
END SDFFNHX2MTH

MACRO SDFFNHX4MTH
    CLASS CORE ;
    FOREIGN SDFFNHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.810 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.078 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 0.990 5.545 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.895 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.1313 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.500 0.765 16.710 1.980 ;
        RECT  16.425 0.765 16.500 1.025 ;
        RECT  16.475 1.720 16.500 1.980 ;
        END
        AntennaDiffArea 0.225 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.595 1.685 15.665 1.945 ;
        RECT  15.335 0.385 15.595 1.945 ;
        RECT  14.820 1.290 15.335 1.580 ;
        RECT  14.530 1.290 14.820 1.945 ;
        END
        AntennaDiffArea 0.762 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.630 1.570 ;
        END
        AntennaGateArea 0.1482 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.240 0.430 1.710 ;
        END
        AntennaGateArea 0.1703 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.105 -0.130 16.810 0.130 ;
        RECT  15.845 -0.130 16.105 0.990 ;
        RECT  15.055 -0.130 15.845 0.130 ;
        RECT  14.455 -0.130 15.055 0.385 ;
        RECT  14.200 -0.130 14.455 0.130 ;
        RECT  13.940 -0.130 14.200 0.515 ;
        RECT  10.330 -0.130 13.940 0.130 ;
        RECT  10.070 -0.130 10.330 0.300 ;
        RECT  8.490 -0.130 10.070 0.130 ;
        RECT  8.230 -0.130 8.490 0.975 ;
        RECT  0.430 -0.130 8.230 0.130 ;
        RECT  0.170 -0.130 0.430 0.300 ;
        RECT  0.000 -0.130 0.170 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.545 2.740 16.810 3.000 ;
        RECT  15.945 2.465 16.545 3.000 ;
        RECT  14.010 2.740 15.945 3.000 ;
        RECT  13.850 1.865 14.010 3.000 ;
        RECT  10.330 2.740 13.850 3.000 ;
        RECT  10.070 2.585 10.330 3.000 ;
        RECT  9.250 2.740 10.070 3.000 ;
        RECT  8.990 2.585 9.250 3.000 ;
        RECT  7.070 2.740 8.990 3.000 ;
        RECT  6.810 2.220 7.070 3.000 ;
        RECT  2.695 2.740 6.810 3.000 ;
        RECT  2.535 2.095 2.695 3.000 ;
        RECT  0.770 2.740 2.535 3.000 ;
        RECT  0.265 2.460 0.770 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.135 1.265 16.295 2.285 ;
        RECT  14.670 2.125 16.135 2.285 ;
        RECT  14.350 0.815 14.670 0.975 ;
        RECT  14.410 2.125 14.670 2.540 ;
        RECT  14.350 2.125 14.410 2.285 ;
        RECT  14.190 0.815 14.350 2.285 ;
        RECT  13.780 1.220 14.190 1.480 ;
        RECT  13.440 0.310 13.600 1.735 ;
        RECT  11.390 0.310 13.440 0.470 ;
        RECT  13.160 1.475 13.440 1.735 ;
        RECT  13.100 0.765 13.260 1.280 ;
        RECT  13.060 1.915 13.170 2.075 ;
        RECT  12.980 1.120 13.100 1.280 ;
        RECT  12.980 1.915 13.060 2.480 ;
        RECT  12.820 1.120 12.980 2.480 ;
        RECT  12.290 1.120 12.820 1.280 ;
        RECT  11.790 2.320 12.820 2.480 ;
        RECT  12.540 0.650 12.800 0.940 ;
        RECT  11.730 0.650 12.540 0.810 ;
        RECT  12.250 1.980 12.350 2.140 ;
        RECT  12.030 0.990 12.290 1.280 ;
        RECT  12.090 1.570 12.250 2.140 ;
        RECT  11.790 1.570 12.090 1.730 ;
        RECT  11.730 1.100 11.790 1.730 ;
        RECT  11.630 2.220 11.790 2.480 ;
        RECT  11.630 0.650 11.730 1.730 ;
        RECT  11.570 0.650 11.630 1.275 ;
        RECT  11.110 1.100 11.570 1.275 ;
        RECT  11.290 1.555 11.450 2.475 ;
        RECT  11.230 0.310 11.390 0.640 ;
        RECT  10.670 2.315 11.290 2.475 ;
        RECT  9.640 0.480 11.230 0.640 ;
        RECT  10.950 0.820 11.110 2.135 ;
        RECT  10.610 0.820 10.950 0.980 ;
        RECT  10.850 1.905 10.950 2.135 ;
        RECT  9.530 1.905 10.850 2.065 ;
        RECT  10.390 1.265 10.730 1.525 ;
        RECT  10.510 2.245 10.670 2.475 ;
        RECT  8.635 2.245 10.510 2.405 ;
        RECT  10.230 0.865 10.390 1.525 ;
        RECT  9.170 0.865 10.230 1.025 ;
        RECT  9.380 0.345 9.640 0.640 ;
        RECT  9.370 1.340 9.530 2.065 ;
        RECT  8.830 0.480 9.380 0.640 ;
        RECT  9.010 0.865 9.170 1.655 ;
        RECT  8.390 1.495 9.010 1.655 ;
        RECT  8.670 0.480 8.830 1.315 ;
        RECT  8.010 1.155 8.670 1.315 ;
        RECT  8.475 2.245 8.635 2.445 ;
        RECT  7.435 2.285 8.475 2.445 ;
        RECT  7.790 1.495 8.390 2.085 ;
        RECT  7.850 0.465 8.010 1.315 ;
        RECT  7.100 0.465 7.850 0.625 ;
        RECT  7.670 1.495 7.790 1.655 ;
        RECT  7.510 0.805 7.670 1.655 ;
        RECT  7.280 0.805 7.510 0.965 ;
        RECT  7.330 1.880 7.435 2.445 ;
        RECT  7.275 1.145 7.330 2.445 ;
        RECT  7.170 1.145 7.275 2.040 ;
        RECT  6.925 1.145 7.170 1.305 ;
        RECT  6.630 1.880 7.170 2.040 ;
        RECT  6.940 0.465 7.100 0.810 ;
        RECT  6.485 1.540 6.990 1.700 ;
        RECT  6.485 0.650 6.940 0.810 ;
        RECT  6.665 0.990 6.925 1.305 ;
        RECT  6.145 0.310 6.760 0.470 ;
        RECT  6.470 1.880 6.630 2.280 ;
        RECT  6.325 0.650 6.485 1.700 ;
        RECT  6.290 2.120 6.470 2.280 ;
        RECT  6.290 1.540 6.325 1.700 ;
        RECT  6.130 1.540 6.290 1.940 ;
        RECT  6.130 2.120 6.290 2.560 ;
        RECT  5.985 0.310 6.145 0.810 ;
        RECT  5.950 1.780 6.130 1.940 ;
        RECT  3.035 2.400 6.130 2.560 ;
        RECT  5.950 0.650 5.985 0.810 ;
        RECT  5.790 0.650 5.950 1.600 ;
        RECT  5.790 1.780 5.950 2.220 ;
        RECT  0.770 0.310 5.805 0.470 ;
        RECT  4.120 0.650 5.790 0.810 ;
        RECT  5.610 1.440 5.790 1.600 ;
        RECT  3.375 2.060 5.790 2.220 ;
        RECT  5.450 1.440 5.610 1.880 ;
        RECT  4.065 1.720 5.450 1.880 ;
        RECT  3.715 1.720 3.815 1.880 ;
        RECT  3.715 0.650 3.750 0.810 ;
        RECT  3.555 0.650 3.715 1.880 ;
        RECT  3.490 0.650 3.555 0.810 ;
        RECT  3.215 1.410 3.375 2.220 ;
        RECT  3.150 0.650 3.310 1.230 ;
        RECT  2.970 1.410 3.215 1.570 ;
        RECT  1.110 0.650 3.150 0.810 ;
        RECT  2.875 1.750 3.035 2.560 ;
        RECT  2.810 0.990 2.970 1.570 ;
        RECT  1.980 1.750 2.875 1.910 ;
        RECT  1.450 0.990 2.810 1.150 ;
        RECT  1.965 2.095 2.125 2.560 ;
        RECT  1.820 1.720 1.980 1.910 ;
        RECT  1.110 2.400 1.965 2.560 ;
        RECT  1.790 1.720 1.820 1.880 ;
        RECT  1.630 1.540 1.790 1.880 ;
        RECT  1.450 2.060 1.665 2.220 ;
        RECT  1.290 0.990 1.450 2.220 ;
        RECT  0.950 0.650 1.110 2.560 ;
        RECT  0.610 0.310 0.770 2.070 ;
        RECT  0.125 0.765 0.610 1.025 ;
        RECT  0.385 1.910 0.610 2.070 ;
        RECT  0.125 1.910 0.385 2.170 ;
    END
END SDFFNHX4MTH

MACRO SDFFNHX8MTH
    CLASS CORE ;
    FOREIGN SDFFNHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.630 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.630 1.330 5.270 1.540 ;
        END
        AntennaGateArea 0.1105 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.370 0.990 5.630 1.180 ;
        RECT  4.450 0.990 5.370 1.150 ;
        RECT  4.290 0.990 4.450 1.540 ;
        RECT  3.945 1.280 4.290 1.540 ;
        END
        AntennaGateArea 0.1651 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.365 0.805 14.660 2.505 ;
        END
        AntennaDiffArea 0.294 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.735 0.385 16.995 2.395 ;
        RECT  16.045 1.330 16.735 1.590 ;
        RECT  16.040 0.385 16.045 1.590 ;
        RECT  15.780 0.385 16.040 2.395 ;
        END
        AntennaDiffArea 1.198 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.630 1.570 ;
        END
        AntennaGateArea 0.1612 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.240 0.430 1.710 ;
        END
        AntennaGateArea 0.2639 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.505 -0.130 17.630 0.130 ;
        RECT  17.245 -0.130 17.505 0.985 ;
        RECT  14.380 -0.130 17.245 0.130 ;
        RECT  13.780 -0.130 14.380 0.280 ;
        RECT  10.330 -0.130 13.780 0.130 ;
        RECT  10.070 -0.130 10.330 0.300 ;
        RECT  8.490 -0.130 10.070 0.130 ;
        RECT  8.230 -0.130 8.490 0.975 ;
        RECT  0.430 -0.130 8.230 0.130 ;
        RECT  0.170 -0.130 0.430 0.300 ;
        RECT  0.000 -0.130 0.170 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.505 2.740 17.630 3.000 ;
        RECT  17.245 1.795 17.505 3.000 ;
        RECT  15.530 2.740 17.245 3.000 ;
        RECT  15.270 2.175 15.530 3.000 ;
        RECT  14.060 2.740 15.270 3.000 ;
        RECT  13.800 1.865 14.060 3.000 ;
        RECT  10.330 2.740 13.800 3.000 ;
        RECT  10.070 2.585 10.330 3.000 ;
        RECT  9.250 2.740 10.070 3.000 ;
        RECT  8.990 2.585 9.250 3.000 ;
        RECT  7.090 2.740 8.990 3.000 ;
        RECT  6.830 2.220 7.090 3.000 ;
        RECT  2.695 2.740 6.830 3.000 ;
        RECT  2.535 2.095 2.695 3.000 ;
        RECT  0.000 2.740 2.535 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.915 0.310 15.075 1.935 ;
        RECT  14.815 0.310 14.915 0.625 ;
        RECT  14.860 1.675 14.915 1.935 ;
        RECT  13.995 0.465 14.815 0.625 ;
        RECT  13.995 1.285 14.095 1.545 ;
        RECT  13.835 0.465 13.995 1.545 ;
        RECT  13.440 0.310 13.600 1.735 ;
        RECT  11.180 0.310 13.440 0.470 ;
        RECT  13.160 1.475 13.440 1.735 ;
        RECT  13.100 0.755 13.260 1.280 ;
        RECT  13.060 1.915 13.170 2.075 ;
        RECT  12.980 1.120 13.100 1.280 ;
        RECT  12.980 1.915 13.060 2.480 ;
        RECT  12.820 1.120 12.980 2.480 ;
        RECT  12.290 1.120 12.820 1.280 ;
        RECT  11.790 2.320 12.820 2.480 ;
        RECT  12.540 0.650 12.800 0.940 ;
        RECT  11.780 0.650 12.540 0.810 ;
        RECT  12.190 1.980 12.350 2.140 ;
        RECT  12.030 0.990 12.290 1.280 ;
        RECT  12.030 1.500 12.190 2.140 ;
        RECT  11.845 1.500 12.030 1.660 ;
        RECT  11.780 1.115 11.845 1.660 ;
        RECT  11.630 1.880 11.790 2.480 ;
        RECT  11.685 0.650 11.780 1.660 ;
        RECT  11.520 0.650 11.685 1.275 ;
        RECT  11.110 1.115 11.520 1.275 ;
        RECT  11.290 1.485 11.450 2.475 ;
        RECT  10.670 2.315 11.290 2.475 ;
        RECT  11.020 0.310 11.180 0.640 ;
        RECT  10.950 0.820 11.110 2.135 ;
        RECT  9.700 0.480 11.020 0.640 ;
        RECT  10.610 0.820 10.950 0.980 ;
        RECT  10.850 1.905 10.950 2.135 ;
        RECT  9.530 1.905 10.850 2.065 ;
        RECT  10.510 2.245 10.670 2.475 ;
        RECT  8.635 2.245 10.510 2.405 ;
        RECT  10.390 1.265 10.500 1.525 ;
        RECT  10.230 0.865 10.390 1.525 ;
        RECT  9.170 0.865 10.230 1.025 ;
        RECT  9.440 0.345 9.700 0.640 ;
        RECT  9.370 1.340 9.530 2.065 ;
        RECT  8.830 0.480 9.440 0.640 ;
        RECT  9.010 0.865 9.170 1.655 ;
        RECT  8.390 1.495 9.010 1.655 ;
        RECT  8.670 0.480 8.830 1.315 ;
        RECT  8.010 1.155 8.670 1.315 ;
        RECT  8.475 2.245 8.635 2.455 ;
        RECT  7.435 2.295 8.475 2.455 ;
        RECT  7.790 1.495 8.390 2.085 ;
        RECT  7.850 0.465 8.010 1.315 ;
        RECT  7.100 0.465 7.850 0.625 ;
        RECT  7.670 1.495 7.790 1.655 ;
        RECT  7.510 0.805 7.670 1.655 ;
        RECT  7.280 0.805 7.510 0.965 ;
        RECT  7.330 1.880 7.435 2.455 ;
        RECT  7.275 1.145 7.330 2.455 ;
        RECT  7.170 1.145 7.275 2.040 ;
        RECT  6.925 1.145 7.170 1.305 ;
        RECT  6.650 1.880 7.170 2.040 ;
        RECT  6.940 0.465 7.100 0.810 ;
        RECT  6.485 1.540 6.990 1.700 ;
        RECT  6.485 0.650 6.940 0.810 ;
        RECT  6.665 0.990 6.925 1.305 ;
        RECT  6.145 0.310 6.760 0.470 ;
        RECT  6.490 1.880 6.650 2.280 ;
        RECT  6.290 2.120 6.490 2.280 ;
        RECT  6.325 0.650 6.485 1.700 ;
        RECT  6.310 1.540 6.325 1.700 ;
        RECT  6.150 1.540 6.310 1.940 ;
        RECT  6.130 2.120 6.290 2.560 ;
        RECT  5.950 1.780 6.150 1.940 ;
        RECT  5.985 0.310 6.145 0.810 ;
        RECT  3.035 2.400 6.130 2.560 ;
        RECT  5.970 0.650 5.985 0.810 ;
        RECT  5.810 0.650 5.970 1.600 ;
        RECT  5.790 1.780 5.950 2.220 ;
        RECT  4.050 0.650 5.810 0.810 ;
        RECT  5.610 1.440 5.810 1.600 ;
        RECT  0.770 0.310 5.805 0.470 ;
        RECT  3.375 2.060 5.790 2.220 ;
        RECT  5.450 1.440 5.610 1.880 ;
        RECT  4.065 1.720 5.450 1.880 ;
        RECT  3.765 1.720 3.815 1.880 ;
        RECT  3.605 0.650 3.765 1.880 ;
        RECT  3.490 0.650 3.605 0.810 ;
        RECT  3.555 1.720 3.605 1.880 ;
        RECT  3.310 0.970 3.405 1.230 ;
        RECT  3.215 1.410 3.375 2.220 ;
        RECT  3.150 0.650 3.310 1.230 ;
        RECT  2.970 1.410 3.215 1.570 ;
        RECT  1.110 0.650 3.150 0.810 ;
        RECT  2.875 1.750 3.035 2.560 ;
        RECT  2.810 0.990 2.970 1.570 ;
        RECT  1.980 1.750 2.875 1.910 ;
        RECT  1.450 0.990 2.810 1.150 ;
        RECT  1.965 2.095 2.125 2.560 ;
        RECT  1.820 1.720 1.980 1.910 ;
        RECT  1.110 2.400 1.965 2.560 ;
        RECT  1.790 1.720 1.820 1.880 ;
        RECT  1.630 1.540 1.790 1.880 ;
        RECT  1.450 2.060 1.665 2.220 ;
        RECT  1.290 0.990 1.450 2.220 ;
        RECT  0.950 0.650 1.110 2.560 ;
        RECT  0.610 0.310 0.770 2.270 ;
        RECT  0.125 0.685 0.610 0.945 ;
        RECT  0.125 2.010 0.610 2.270 ;
    END
END SDFFNHX8MTH

MACRO SDFFNSRHX1MTH
    CLASS CORE ;
    FOREIGN SDFFNSRHX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.220 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 1.145 6.935 1.660 ;
        END
        AntennaGateArea 0.1391 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.935 1.330 4.260 1.540 ;
        RECT  3.775 1.330 3.935 1.715 ;
        RECT  3.750 1.330 3.775 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.990 4.775 1.150 ;
        RECT  3.540 1.700 3.590 1.990 ;
        RECT  3.380 0.990 3.540 1.990 ;
        RECT  3.195 0.990 3.380 1.475 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.080 1.385 13.315 1.545 ;
        RECT  11.920 1.385 12.080 1.635 ;
        RECT  11.010 1.475 11.920 1.635 ;
        RECT  10.530 1.330 11.010 1.635 ;
        END
        AntennaGateArea 0.1417 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.480 2.245 15.965 2.405 ;
        RECT  15.210 2.065 15.480 2.405 ;
        RECT  15.210 0.815 15.425 0.975 ;
        RECT  15.050 0.815 15.210 2.405 ;
        END
        AntennaDiffArea 0.342 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.885 0.765 17.120 2.285 ;
        END
        AntennaDiffArea 0.34 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.255 2.675 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.225 0.895 1.580 ;
        END
        AntennaGateArea 0.1469 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.675 -0.130 17.220 0.130 ;
        RECT  15.735 -0.130 16.675 0.260 ;
        RECT  2.335 -0.130 15.735 0.130 ;
        RECT  1.735 -0.130 2.335 0.250 ;
        RECT  0.810 -0.130 1.735 0.130 ;
        RECT  0.210 -0.130 0.810 0.250 ;
        RECT  0.000 -0.130 0.210 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.585 2.740 17.220 3.000 ;
        RECT  16.325 1.685 16.585 3.000 ;
        RECT  11.505 2.740 16.325 3.000 ;
        RECT  10.905 2.620 11.505 3.000 ;
        RECT  10.110 2.740 10.905 3.000 ;
        RECT  9.850 2.620 10.110 3.000 ;
        RECT  9.085 2.740 9.850 3.000 ;
        RECT  8.485 2.620 9.085 3.000 ;
        RECT  6.865 2.740 8.485 3.000 ;
        RECT  6.265 2.620 6.865 3.000 ;
        RECT  2.635 2.740 6.265 3.000 ;
        RECT  2.375 2.620 2.635 3.000 ;
        RECT  0.755 2.740 2.375 3.000 ;
        RECT  0.255 2.365 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.535 1.185 16.705 1.445 ;
        RECT  16.375 0.475 16.535 1.445 ;
        RECT  14.870 0.475 16.375 0.635 ;
        RECT  16.205 1.185 16.375 1.445 ;
        RECT  15.965 0.815 16.125 0.975 ;
        RECT  15.805 0.815 15.965 1.945 ;
        RECT  15.415 1.240 15.805 1.840 ;
        RECT  14.710 0.355 14.870 2.505 ;
        RECT  14.305 0.355 14.710 0.550 ;
        RECT  14.110 2.295 14.710 2.505 ;
        RECT  14.490 1.500 14.530 1.760 ;
        RECT  14.390 0.760 14.490 1.760 ;
        RECT  14.230 0.760 14.390 2.115 ;
        RECT  12.430 0.355 14.305 0.515 ;
        RECT  13.655 1.955 14.230 2.115 ;
        RECT  12.820 2.295 14.110 2.455 ;
        RECT  13.890 0.695 14.050 1.775 ;
        RECT  12.250 0.695 13.890 0.855 ;
        RECT  13.495 1.035 13.655 2.115 ;
        RECT  11.910 1.035 13.495 1.195 ;
        RECT  13.050 1.865 13.495 2.115 ;
        RECT  12.310 2.185 12.635 2.440 ;
        RECT  11.780 1.815 12.540 1.975 ;
        RECT  9.520 2.280 12.310 2.440 ;
        RECT  12.090 0.310 12.250 0.855 ;
        RECT  2.675 0.310 12.090 0.470 ;
        RECT  11.750 0.650 11.910 1.195 ;
        RECT  11.620 1.815 11.780 2.100 ;
        RECT  6.480 0.650 11.750 0.810 ;
        RECT  9.950 1.940 11.620 2.100 ;
        RECT  11.410 0.990 11.570 1.250 ;
        RECT  9.950 0.990 11.410 1.150 ;
        RECT  9.790 0.990 9.950 2.100 ;
        RECT  9.450 0.990 9.610 2.100 ;
        RECT  9.260 2.280 9.520 2.470 ;
        RECT  8.470 1.910 9.450 2.100 ;
        RECT  8.305 2.280 9.260 2.440 ;
        RECT  8.310 0.990 8.470 2.100 ;
        RECT  8.145 0.990 8.310 1.150 ;
        RECT  7.965 1.860 8.310 2.100 ;
        RECT  8.135 2.280 8.305 2.480 ;
        RECT  7.620 2.320 8.135 2.480 ;
        RECT  7.960 1.335 8.100 1.595 ;
        RECT  7.805 1.860 7.965 2.130 ;
        RECT  7.800 1.130 7.960 1.595 ;
        RECT  7.280 1.130 7.800 1.290 ;
        RECT  7.460 1.470 7.620 2.480 ;
        RECT  7.450 2.280 7.460 2.480 ;
        RECT  6.075 2.280 7.450 2.440 ;
        RECT  7.120 1.130 7.280 2.100 ;
        RECT  6.040 1.940 7.120 2.100 ;
        RECT  6.220 0.650 6.480 1.760 ;
        RECT  5.915 2.280 6.075 2.560 ;
        RECT  5.880 0.650 6.040 2.100 ;
        RECT  3.045 2.400 5.915 2.560 ;
        RECT  5.115 0.650 5.880 0.810 ;
        RECT  5.540 0.990 5.700 2.220 ;
        RECT  5.300 0.990 5.540 1.150 ;
        RECT  5.060 2.060 5.540 2.220 ;
        RECT  4.955 0.650 5.115 1.490 ;
        RECT  4.800 1.670 5.060 2.220 ;
        RECT  3.825 0.650 4.955 0.810 ;
        RECT  4.620 1.330 4.955 1.490 ;
        RECT  3.935 2.060 4.800 2.220 ;
        RECT  4.460 1.330 4.620 1.880 ;
        RECT  4.115 1.720 4.460 1.880 ;
        RECT  3.775 1.895 3.935 2.220 ;
        RECT  3.015 0.650 3.515 0.810 ;
        RECT  3.015 1.835 3.155 2.095 ;
        RECT  2.855 2.280 3.045 2.560 ;
        RECT  2.855 0.650 3.015 2.095 ;
        RECT  2.025 2.280 2.855 2.440 ;
        RECT  2.515 0.310 2.675 0.590 ;
        RECT  1.605 0.430 2.515 0.590 ;
        RECT  1.965 0.815 2.045 0.975 ;
        RECT  1.965 2.215 2.025 2.475 ;
        RECT  1.785 0.815 1.965 2.475 ;
        RECT  1.595 1.400 1.785 1.560 ;
        RECT  1.445 0.430 1.605 1.010 ;
        RECT  1.415 1.740 1.605 2.000 ;
        RECT  1.415 0.850 1.445 1.010 ;
        RECT  1.205 0.850 1.415 2.000 ;
        RECT  1.005 0.310 1.265 0.670 ;
        RECT  0.385 0.490 1.005 0.670 ;
        RECT  0.330 0.490 0.385 1.025 ;
        RECT  0.330 1.740 0.360 2.000 ;
        RECT  0.125 0.490 0.330 2.000 ;
    END
END SDFFNSRHX1MTH

MACRO SDFFNSRHX2MTH
    CLASS CORE ;
    FOREIGN SDFFNSRHX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.220 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 1.145 6.935 1.660 ;
        END
        AntennaGateArea 0.1625 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.935 1.330 4.260 1.540 ;
        RECT  3.775 1.330 3.935 1.715 ;
        RECT  3.750 1.330 3.775 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.990 4.775 1.150 ;
        RECT  3.540 1.700 3.590 1.990 ;
        RECT  3.380 0.990 3.540 1.990 ;
        RECT  3.195 0.990 3.380 1.475 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.910 1.385 13.315 1.545 ;
        RECT  11.750 1.385 11.910 1.635 ;
        RECT  11.010 1.475 11.750 1.635 ;
        RECT  10.580 1.330 11.010 1.635 ;
        END
        AntennaGateArea 0.1716 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.480 2.255 15.965 2.415 ;
        RECT  15.235 2.065 15.480 2.415 ;
        RECT  15.235 0.815 15.335 0.975 ;
        RECT  15.075 0.815 15.235 2.415 ;
        END
        AntennaDiffArea 0.401 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.885 0.400 17.120 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.145 1.255 2.675 1.580 ;
        END
        AntennaGateArea 0.0884 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.225 1.000 1.580 ;
        END
        AntennaGateArea 0.1469 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.430 -0.130 17.220 0.130 ;
        RECT  15.830 -0.130 16.430 0.260 ;
        RECT  2.335 -0.130 15.830 0.130 ;
        RECT  1.735 -0.130 2.335 0.250 ;
        RECT  0.810 -0.130 1.735 0.130 ;
        RECT  0.210 -0.130 0.810 0.250 ;
        RECT  0.000 -0.130 0.210 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.585 2.740 17.220 3.000 ;
        RECT  16.325 1.830 16.585 3.000 ;
        RECT  11.100 2.740 16.325 3.000 ;
        RECT  10.840 2.620 11.100 3.000 ;
        RECT  10.160 2.740 10.840 3.000 ;
        RECT  9.900 2.620 10.160 3.000 ;
        RECT  9.010 2.740 9.900 3.000 ;
        RECT  8.750 2.620 9.010 3.000 ;
        RECT  7.420 2.740 8.750 3.000 ;
        RECT  7.160 2.620 7.420 3.000 ;
        RECT  6.820 2.740 7.160 3.000 ;
        RECT  6.220 2.620 6.820 3.000 ;
        RECT  2.640 2.740 6.220 3.000 ;
        RECT  2.380 2.575 2.640 3.000 ;
        RECT  0.805 2.740 2.380 3.000 ;
        RECT  0.205 2.290 0.805 3.000 ;
        RECT  0.000 2.740 0.205 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.535 1.185 16.695 1.445 ;
        RECT  16.375 0.475 16.535 1.445 ;
        RECT  14.870 0.475 16.375 0.635 ;
        RECT  16.195 1.185 16.375 1.445 ;
        RECT  15.965 0.815 15.995 0.975 ;
        RECT  15.805 0.815 15.965 1.945 ;
        RECT  15.735 0.815 15.805 1.840 ;
        RECT  15.415 1.240 15.735 1.840 ;
        RECT  14.710 0.355 14.870 2.505 ;
        RECT  14.305 0.355 14.710 0.550 ;
        RECT  14.110 2.295 14.710 2.505 ;
        RECT  14.370 0.760 14.530 2.115 ;
        RECT  14.230 0.760 14.370 0.920 ;
        RECT  13.655 1.955 14.370 2.115 ;
        RECT  12.430 0.355 14.305 0.515 ;
        RECT  12.820 2.295 14.110 2.455 ;
        RECT  13.890 0.695 14.050 1.775 ;
        RECT  12.250 0.695 13.890 0.855 ;
        RECT  13.495 1.035 13.655 2.115 ;
        RECT  11.910 1.035 13.495 1.195 ;
        RECT  13.050 1.865 13.495 2.115 ;
        RECT  11.780 1.815 12.540 1.975 ;
        RECT  11.995 2.185 12.255 2.440 ;
        RECT  12.090 0.310 12.250 0.855 ;
        RECT  2.675 0.310 12.090 0.470 ;
        RECT  9.570 2.270 11.995 2.440 ;
        RECT  11.750 0.650 11.910 1.195 ;
        RECT  11.620 1.815 11.780 2.090 ;
        RECT  6.480 0.650 11.750 0.810 ;
        RECT  10.000 1.930 11.620 2.090 ;
        RECT  11.410 0.990 11.570 1.250 ;
        RECT  10.000 0.990 11.410 1.150 ;
        RECT  9.840 0.990 10.000 2.090 ;
        RECT  9.310 2.270 9.570 2.560 ;
        RECT  9.400 1.025 9.560 2.090 ;
        RECT  9.110 1.840 9.400 2.090 ;
        RECT  8.440 2.270 9.310 2.440 ;
        RECT  8.610 1.840 9.110 2.000 ;
        RECT  8.450 0.990 8.610 2.000 ;
        RECT  8.260 0.990 8.450 1.150 ;
        RECT  8.100 1.840 8.450 2.000 ;
        RECT  8.280 2.270 8.440 2.480 ;
        RECT  7.740 2.300 8.280 2.480 ;
        RECT  8.080 1.335 8.270 1.595 ;
        RECT  7.940 1.840 8.100 2.120 ;
        RECT  7.920 1.130 8.080 1.595 ;
        RECT  7.400 1.130 7.920 1.290 ;
        RECT  7.600 1.470 7.740 2.480 ;
        RECT  7.580 1.470 7.600 2.440 ;
        RECT  6.040 2.280 7.580 2.440 ;
        RECT  7.240 1.130 7.400 2.100 ;
        RECT  6.040 1.940 7.240 2.100 ;
        RECT  6.220 0.650 6.480 1.760 ;
        RECT  5.880 0.650 6.040 2.100 ;
        RECT  5.880 2.280 6.040 2.560 ;
        RECT  5.115 0.650 5.880 0.810 ;
        RECT  3.140 2.400 5.880 2.560 ;
        RECT  5.540 0.990 5.700 2.220 ;
        RECT  5.300 0.990 5.540 1.150 ;
        RECT  5.060 2.060 5.540 2.220 ;
        RECT  4.955 0.650 5.115 1.490 ;
        RECT  4.800 1.670 5.060 2.220 ;
        RECT  3.825 0.650 4.955 0.810 ;
        RECT  4.620 1.330 4.955 1.490 ;
        RECT  3.935 2.060 4.800 2.220 ;
        RECT  4.460 1.330 4.620 1.880 ;
        RECT  4.115 1.720 4.460 1.880 ;
        RECT  3.775 1.895 3.935 2.220 ;
        RECT  3.015 0.650 3.515 0.810 ;
        RECT  3.015 1.690 3.155 1.950 ;
        RECT  2.955 2.225 3.140 2.560 ;
        RECT  2.855 0.650 3.015 1.950 ;
        RECT  2.110 2.225 2.955 2.390 ;
        RECT  2.515 0.310 2.675 0.635 ;
        RECT  1.605 0.475 2.515 0.635 ;
        RECT  1.965 2.225 2.110 2.485 ;
        RECT  1.965 0.815 2.075 0.975 ;
        RECT  1.785 0.815 1.965 2.485 ;
        RECT  1.535 1.300 1.785 1.560 ;
        RECT  1.445 0.475 1.605 1.010 ;
        RECT  1.355 1.740 1.605 2.000 ;
        RECT  1.355 0.850 1.445 1.010 ;
        RECT  1.195 0.850 1.355 2.000 ;
        RECT  1.005 0.310 1.265 0.670 ;
        RECT  0.385 0.490 1.005 0.670 ;
        RECT  0.330 0.490 0.385 1.025 ;
        RECT  0.330 1.740 0.385 2.000 ;
        RECT  0.125 0.490 0.330 2.000 ;
    END
END SDFFNSRHX2MTH

MACRO SDFFNSRHX4MTH
    CLASS CORE ;
    FOREIGN SDFFNSRHX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.630 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 1.030 7.025 1.670 ;
        END
        AntennaGateArea 0.182 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.930 1.330 4.260 1.540 ;
        RECT  3.750 1.330 3.930 1.610 ;
        RECT  3.720 1.330 3.750 1.540 ;
        END
        AntennaGateArea 0.078 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.990 4.775 1.150 ;
        RECT  3.540 1.700 3.590 1.990 ;
        RECT  3.380 0.990 3.540 1.990 ;
        RECT  3.195 0.990 3.380 1.405 ;
        END
        AntennaGateArea 0.13 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.910 1.385 13.315 1.545 ;
        RECT  11.750 1.385 11.910 1.635 ;
        RECT  11.010 1.475 11.750 1.635 ;
        RECT  10.580 1.330 11.010 1.635 ;
        END
        AntennaGateArea 0.2093 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.480 2.255 15.965 2.415 ;
        RECT  15.235 2.065 15.480 2.415 ;
        RECT  15.235 0.815 15.405 0.975 ;
        RECT  15.075 0.815 15.235 2.415 ;
        END
        AntennaDiffArea 0.351 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.105 1.290 17.195 1.580 ;
        RECT  16.910 0.400 17.105 2.285 ;
        RECT  16.775 0.400 16.910 1.000 ;
        RECT  16.775 1.685 16.910 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.365 1.150 2.675 1.410 ;
        RECT  2.145 1.150 2.365 1.990 ;
        END
        AntennaGateArea 0.156 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.225 0.895 1.580 ;
        END
        AntennaGateArea 0.1664 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.445 -0.130 17.630 0.130 ;
        RECT  17.285 -0.130 17.445 1.000 ;
        RECT  16.390 -0.130 17.285 0.130 ;
        RECT  15.790 -0.130 16.390 0.260 ;
        RECT  0.785 -0.130 15.790 0.130 ;
        RECT  0.185 -0.130 0.785 0.250 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.445 2.740 17.630 3.000 ;
        RECT  17.285 1.815 17.445 3.000 ;
        RECT  16.475 2.740 17.285 3.000 ;
        RECT  16.215 2.255 16.475 3.000 ;
        RECT  10.145 2.740 16.215 3.000 ;
        RECT  9.885 2.620 10.145 3.000 ;
        RECT  8.985 2.740 9.885 3.000 ;
        RECT  8.725 2.620 8.985 3.000 ;
        RECT  6.910 2.740 8.725 3.000 ;
        RECT  6.310 2.620 6.910 3.000 ;
        RECT  2.640 2.740 6.310 3.000 ;
        RECT  2.380 2.575 2.640 3.000 ;
        RECT  0.755 2.740 2.380 3.000 ;
        RECT  0.255 2.365 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.535 1.185 16.695 1.445 ;
        RECT  16.375 0.475 16.535 1.445 ;
        RECT  14.870 0.475 16.375 0.635 ;
        RECT  16.195 1.185 16.375 1.445 ;
        RECT  15.965 0.815 16.015 0.975 ;
        RECT  15.755 0.815 15.965 1.945 ;
        RECT  15.415 1.240 15.755 1.840 ;
        RECT  14.710 0.355 14.870 2.505 ;
        RECT  14.470 0.355 14.710 0.550 ;
        RECT  14.110 2.295 14.710 2.505 ;
        RECT  14.370 0.760 14.530 2.115 ;
        RECT  12.430 0.355 14.470 0.515 ;
        RECT  14.270 0.760 14.370 0.920 ;
        RECT  13.655 1.955 14.370 2.115 ;
        RECT  12.820 2.295 14.110 2.455 ;
        RECT  13.890 0.695 14.050 1.775 ;
        RECT  12.250 0.695 13.890 0.855 ;
        RECT  13.495 1.035 13.655 2.115 ;
        RECT  11.910 1.035 13.495 1.195 ;
        RECT  13.050 1.865 13.495 2.115 ;
        RECT  11.780 1.815 12.540 1.975 ;
        RECT  11.995 2.185 12.255 2.440 ;
        RECT  12.090 0.310 12.250 0.855 ;
        RECT  1.605 0.310 12.090 0.470 ;
        RECT  9.570 2.270 11.995 2.440 ;
        RECT  11.750 0.650 11.910 1.195 ;
        RECT  11.620 1.815 11.780 2.090 ;
        RECT  6.480 0.650 11.750 0.810 ;
        RECT  9.985 1.930 11.620 2.090 ;
        RECT  11.410 0.990 11.570 1.250 ;
        RECT  9.985 0.990 11.410 1.150 ;
        RECT  9.825 0.990 9.985 2.090 ;
        RECT  9.295 2.270 9.570 2.560 ;
        RECT  9.400 1.055 9.560 2.090 ;
        RECT  9.095 1.860 9.400 2.090 ;
        RECT  8.440 2.270 9.295 2.440 ;
        RECT  8.610 1.860 9.095 2.020 ;
        RECT  8.450 0.990 8.610 2.020 ;
        RECT  8.260 0.990 8.450 1.150 ;
        RECT  8.100 1.860 8.450 2.020 ;
        RECT  8.280 2.270 8.440 2.470 ;
        RECT  7.740 2.300 8.280 2.470 ;
        RECT  8.080 1.335 8.255 1.595 ;
        RECT  7.925 1.860 8.100 2.120 ;
        RECT  7.920 1.130 8.080 1.595 ;
        RECT  7.400 1.130 7.920 1.290 ;
        RECT  7.600 1.495 7.740 2.470 ;
        RECT  7.580 1.495 7.600 2.440 ;
        RECT  6.075 2.280 7.580 2.440 ;
        RECT  7.240 1.130 7.400 2.100 ;
        RECT  6.040 1.940 7.240 2.100 ;
        RECT  6.220 0.650 6.480 1.760 ;
        RECT  5.915 2.280 6.075 2.560 ;
        RECT  5.880 0.650 6.040 2.100 ;
        RECT  3.140 2.400 5.915 2.560 ;
        RECT  5.115 0.650 5.880 0.810 ;
        RECT  5.540 0.990 5.700 2.220 ;
        RECT  5.300 0.990 5.540 1.150 ;
        RECT  5.060 2.060 5.540 2.220 ;
        RECT  4.955 0.650 5.115 1.490 ;
        RECT  4.800 1.670 5.060 2.220 ;
        RECT  3.825 0.650 4.955 0.810 ;
        RECT  4.620 1.330 4.955 1.490 ;
        RECT  3.935 2.060 4.800 2.220 ;
        RECT  4.460 1.330 4.620 1.880 ;
        RECT  4.115 1.720 4.460 1.880 ;
        RECT  3.775 1.885 3.935 2.220 ;
        RECT  3.015 0.650 3.400 0.810 ;
        RECT  3.015 1.690 3.155 1.950 ;
        RECT  2.955 2.225 3.140 2.560 ;
        RECT  2.855 0.650 3.015 1.950 ;
        RECT  2.150 2.225 2.955 2.390 ;
        RECT  1.965 2.225 2.150 2.525 ;
        RECT  1.965 0.650 2.075 0.810 ;
        RECT  1.785 0.650 1.965 2.525 ;
        RECT  1.575 1.285 1.785 1.545 ;
        RECT  1.445 0.310 1.605 1.010 ;
        RECT  1.320 1.740 1.605 2.000 ;
        RECT  1.320 0.790 1.445 1.010 ;
        RECT  1.095 0.790 1.320 2.000 ;
        RECT  1.005 0.310 1.265 0.610 ;
        RECT  0.385 0.430 1.005 0.610 ;
        RECT  0.310 0.430 0.385 1.025 ;
        RECT  0.310 1.740 0.385 2.000 ;
        RECT  0.125 0.430 0.310 2.000 ;
    END
END SDFFNSRHX4MTH

MACRO SDFFNSRHX8MTH
    CLASS CORE ;
    FOREIGN SDFFNSRHX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 19.270 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.070 1.230 7.460 1.740 ;
        END
        AntennaGateArea 0.2262 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.375 1.330 4.670 1.540 ;
        RECT  4.160 1.330 4.375 1.610 ;
        END
        AntennaGateArea 0.1391 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.950 0.990 5.190 1.150 ;
        RECT  3.950 1.700 4.000 1.990 ;
        RECT  3.790 0.990 3.950 1.990 ;
        RECT  3.635 0.990 3.790 1.475 ;
        END
        AntennaGateArea 0.195 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.320 1.385 13.725 1.545 ;
        RECT  12.160 1.385 12.320 1.635 ;
        RECT  11.420 1.475 12.160 1.635 ;
        RECT  10.990 1.330 11.420 1.635 ;
        END
        AntennaGateArea 0.2119 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.645 2.150 16.545 2.415 ;
        RECT  15.645 0.815 15.815 0.975 ;
        RECT  15.485 0.815 15.645 2.415 ;
        END
        AntennaDiffArea 0.351 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.340 0.400 18.600 2.285 ;
        RECT  17.580 0.905 18.340 1.065 ;
        RECT  17.895 1.330 18.340 1.745 ;
        RECT  17.580 1.585 17.895 1.745 ;
        RECT  17.320 0.400 17.580 1.065 ;
        RECT  17.320 1.585 17.580 2.285 ;
        END
        AntennaDiffArea 1.204 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 0.990 3.115 1.315 ;
        RECT  2.560 0.990 2.770 1.580 ;
        END
        AntennaGateArea 0.2041 ;
    END D
    PIN CKN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.195 0.925 1.580 ;
        END
        AntennaGateArea 0.26 ;
    END CKN
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.110 -0.130 19.270 0.130 ;
        RECT  18.850 -0.130 19.110 1.000 ;
        RECT  18.090 -0.130 18.850 0.130 ;
        RECT  17.830 -0.130 18.090 0.705 ;
        RECT  16.840 -0.130 17.830 0.130 ;
        RECT  16.240 -0.130 16.840 0.260 ;
        RECT  0.775 -0.130 16.240 0.130 ;
        RECT  0.175 -0.130 0.775 0.250 ;
        RECT  0.000 -0.130 0.175 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.110 2.740 19.270 3.000 ;
        RECT  18.850 1.815 19.110 3.000 ;
        RECT  18.090 2.740 18.850 3.000 ;
        RECT  17.830 1.965 18.090 3.000 ;
        RECT  17.070 2.740 17.830 3.000 ;
        RECT  16.810 1.840 17.070 3.000 ;
        RECT  10.570 2.740 16.810 3.000 ;
        RECT  10.310 2.620 10.570 3.000 ;
        RECT  9.420 2.740 10.310 3.000 ;
        RECT  9.160 2.620 9.420 3.000 ;
        RECT  7.355 2.740 9.160 3.000 ;
        RECT  6.755 2.620 7.355 3.000 ;
        RECT  2.005 2.740 6.755 3.000 ;
        RECT  1.805 2.530 2.005 3.000 ;
        RECT  0.735 2.740 1.805 3.000 ;
        RECT  0.235 2.530 0.735 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  17.030 1.245 17.555 1.405 ;
        RECT  16.870 0.475 17.030 1.405 ;
        RECT  15.280 0.475 16.870 0.635 ;
        RECT  16.615 1.245 16.870 1.405 ;
        RECT  16.375 1.685 16.450 1.945 ;
        RECT  16.375 0.815 16.425 0.975 ;
        RECT  16.165 0.815 16.375 1.945 ;
        RECT  15.825 1.240 16.165 1.840 ;
        RECT  15.120 0.355 15.280 2.505 ;
        RECT  14.755 0.355 15.120 0.565 ;
        RECT  14.520 2.295 15.120 2.505 ;
        RECT  14.780 0.775 14.940 2.115 ;
        RECT  14.680 0.775 14.780 0.935 ;
        RECT  14.065 1.955 14.780 2.115 ;
        RECT  12.840 0.355 14.755 0.515 ;
        RECT  13.230 2.295 14.520 2.455 ;
        RECT  14.410 1.615 14.510 1.775 ;
        RECT  14.250 0.695 14.410 1.775 ;
        RECT  12.660 0.695 14.250 0.855 ;
        RECT  13.905 1.035 14.065 2.115 ;
        RECT  12.320 1.035 13.905 1.195 ;
        RECT  13.460 1.865 13.905 2.115 ;
        RECT  12.190 1.815 12.950 1.975 ;
        RECT  12.430 2.185 12.690 2.440 ;
        RECT  12.500 0.310 12.660 0.855 ;
        RECT  1.745 0.310 12.500 0.470 ;
        RECT  9.980 2.270 12.430 2.440 ;
        RECT  12.160 0.650 12.320 1.195 ;
        RECT  12.030 1.815 12.190 2.090 ;
        RECT  6.840 0.650 12.160 0.810 ;
        RECT  10.410 1.930 12.030 2.090 ;
        RECT  11.820 0.990 11.980 1.250 ;
        RECT  10.410 0.990 11.820 1.150 ;
        RECT  10.250 0.990 10.410 2.090 ;
        RECT  9.910 0.990 10.070 2.085 ;
        RECT  9.720 2.270 9.980 2.560 ;
        RECT  9.520 1.860 9.910 2.085 ;
        RECT  8.850 2.270 9.720 2.430 ;
        RECT  9.020 1.860 9.520 2.020 ;
        RECT  8.860 0.990 9.020 2.020 ;
        RECT  8.670 0.990 8.860 1.150 ;
        RECT  8.510 1.860 8.860 2.020 ;
        RECT  8.690 2.270 8.850 2.470 ;
        RECT  8.150 2.300 8.690 2.470 ;
        RECT  8.490 1.335 8.680 1.595 ;
        RECT  8.350 1.860 8.510 2.120 ;
        RECT  8.330 1.130 8.490 1.595 ;
        RECT  7.810 1.130 8.330 1.290 ;
        RECT  8.010 1.495 8.150 2.470 ;
        RECT  7.990 1.495 8.010 2.440 ;
        RECT  6.485 2.280 7.990 2.440 ;
        RECT  7.650 1.130 7.810 2.100 ;
        RECT  6.450 1.940 7.650 2.100 ;
        RECT  6.840 1.600 6.890 1.760 ;
        RECT  6.630 0.650 6.840 1.760 ;
        RECT  6.325 2.280 6.485 2.560 ;
        RECT  6.290 0.650 6.450 2.100 ;
        RECT  2.575 2.400 6.325 2.560 ;
        RECT  5.530 0.650 6.290 0.810 ;
        RECT  5.950 0.990 6.110 2.220 ;
        RECT  5.710 0.990 5.950 1.150 ;
        RECT  5.475 2.060 5.950 2.220 ;
        RECT  5.370 0.650 5.530 1.490 ;
        RECT  5.215 1.670 5.475 2.220 ;
        RECT  4.235 0.650 5.370 0.810 ;
        RECT  5.030 1.330 5.370 1.490 ;
        RECT  4.365 2.060 5.215 2.220 ;
        RECT  4.870 1.330 5.030 1.880 ;
        RECT  4.530 1.720 4.870 1.880 ;
        RECT  4.205 1.960 4.365 2.220 ;
        RECT  3.455 0.650 3.810 0.810 ;
        RECT  3.455 2.060 3.590 2.220 ;
        RECT  3.295 0.650 3.455 2.220 ;
        RECT  2.380 1.870 2.575 2.560 ;
        RECT  2.380 0.650 2.515 0.810 ;
        RECT  2.200 0.650 2.380 2.560 ;
        RECT  1.535 1.285 2.200 1.545 ;
        RECT  1.585 0.310 1.745 1.010 ;
        RECT  1.350 1.740 1.635 2.000 ;
        RECT  1.350 0.790 1.585 1.010 ;
        RECT  1.145 0.790 1.350 2.000 ;
        RECT  1.035 0.310 1.295 0.610 ;
        RECT  0.385 0.430 1.035 0.610 ;
        RECT  0.310 0.430 0.385 1.025 ;
        RECT  0.310 1.835 0.385 2.095 ;
        RECT  0.125 0.430 0.310 2.095 ;
    END
END SDFFNSRHX8MTH

MACRO SDFFQNX1MTH
    CLASS CORE ;
    FOREIGN SDFFQNX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.160 1.950 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.760 2.120 1.920 ;
        RECT  1.130 1.355 1.255 1.920 ;
        RECT  1.095 1.290 1.130 1.920 ;
        RECT  0.915 1.290 1.095 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.165 0.735 9.330 2.115 ;
        RECT  9.045 0.735 9.165 0.995 ;
        RECT  9.055 1.685 9.165 2.115 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.360 1.580 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.700 4.665 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 -0.130 9.430 0.130 ;
        RECT  8.015 -0.130 8.615 0.250 ;
        RECT  6.615 -0.130 8.015 0.130 ;
        RECT  6.065 -0.130 6.615 0.325 ;
        RECT  0.385 -0.130 6.065 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 2.740 9.430 3.000 ;
        RECT  8.110 2.570 8.710 3.000 ;
        RECT  6.530 2.740 8.110 3.000 ;
        RECT  6.270 2.620 6.530 3.000 ;
        RECT  5.645 2.740 6.270 3.000 ;
        RECT  5.045 2.620 5.645 3.000 ;
        RECT  4.250 2.740 5.045 3.000 ;
        RECT  3.990 2.620 4.250 3.000 ;
        RECT  1.920 2.740 3.990 3.000 ;
        RECT  1.660 2.490 1.920 3.000 ;
        RECT  0.000 2.740 1.660 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.875 1.215 8.985 1.475 ;
        RECT  8.715 1.215 8.875 2.105 ;
        RECT  8.095 1.945 8.715 2.105 ;
        RECT  8.375 0.430 8.535 1.405 ;
        RECT  7.755 0.430 8.375 0.590 ;
        RECT  8.345 1.145 8.375 1.405 ;
        RECT  8.095 0.815 8.195 0.975 ;
        RECT  7.935 0.815 8.095 2.105 ;
        RECT  7.830 1.525 7.935 1.785 ;
        RECT  7.595 0.430 7.755 1.300 ;
        RECT  6.915 0.430 7.595 0.590 ;
        RECT  7.530 1.140 7.595 1.300 ;
        RECT  7.370 1.140 7.530 2.465 ;
        RECT  7.190 0.800 7.415 0.960 ;
        RECT  7.150 2.305 7.370 2.465 ;
        RECT  7.030 0.800 7.190 2.105 ;
        RECT  6.965 1.945 7.030 2.105 ;
        RECT  6.805 1.945 6.965 2.440 ;
        RECT  6.690 1.360 6.850 1.620 ;
        RECT  6.085 2.280 6.805 2.440 ;
        RECT  6.220 1.360 6.690 1.520 ;
        RECT  6.365 1.915 6.625 2.100 ;
        RECT  5.665 1.940 6.365 2.100 ;
        RECT  5.960 1.360 6.220 1.760 ;
        RECT  5.825 2.280 6.085 2.540 ;
        RECT  5.890 1.360 5.960 1.520 ;
        RECT  5.755 0.680 5.890 1.520 ;
        RECT  3.795 2.280 5.825 2.440 ;
        RECT  5.730 0.325 5.755 1.520 ;
        RECT  5.595 0.325 5.730 0.840 ;
        RECT  5.505 1.815 5.665 2.100 ;
        RECT  3.160 0.325 5.595 0.485 ;
        RECT  5.295 1.815 5.505 1.975 ;
        RECT  5.135 0.795 5.295 1.975 ;
        RECT  4.980 1.355 5.135 1.975 ;
        RECT  3.880 1.355 4.980 1.515 ;
        RECT  4.765 0.670 4.925 1.165 ;
        RECT  3.435 1.005 4.765 1.165 ;
        RECT  2.960 0.665 4.540 0.825 ;
        RECT  3.635 2.280 3.795 2.560 ;
        RECT  3.385 2.345 3.635 2.560 ;
        RECT  3.275 1.005 3.435 2.165 ;
        RECT  3.095 2.345 3.385 2.505 ;
        RECT  3.140 1.005 3.275 1.195 ;
        RECT  2.925 1.035 3.140 1.195 ;
        RECT  2.935 1.375 3.095 2.505 ;
        RECT  2.800 0.665 2.960 0.855 ;
        RECT  2.745 1.375 2.935 1.535 ;
        RECT  2.745 0.695 2.800 0.855 ;
        RECT  2.595 1.905 2.755 2.505 ;
        RECT  2.585 0.695 2.745 1.535 ;
        RECT  0.660 0.355 2.620 0.515 ;
        RECT  0.970 2.125 2.595 2.285 ;
        RECT  1.665 0.695 1.925 0.890 ;
        RECT  0.915 0.695 1.665 0.855 ;
        RECT  0.810 2.125 0.970 2.505 ;
        RECT  0.655 0.695 0.915 1.075 ;
        RECT  0.630 1.785 0.830 1.945 ;
        RECT  0.630 0.885 0.655 1.075 ;
        RECT  0.350 0.885 0.630 2.560 ;
    END
END SDFFQNX1MTH

MACRO SDFFQNX2MTH
    CLASS CORE ;
    FOREIGN SDFFQNX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.160 1.950 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.760 2.120 1.920 ;
        RECT  1.130 1.355 1.255 1.920 ;
        RECT  1.095 1.290 1.130 1.920 ;
        RECT  0.915 1.290 1.095 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.165 0.425 9.330 2.285 ;
        RECT  9.045 0.425 9.165 1.025 ;
        RECT  9.075 1.685 9.165 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.360 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.695 4.665 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.615 -0.130 9.430 0.130 ;
        RECT  8.015 -0.130 8.615 0.250 ;
        RECT  6.615 -0.130 8.015 0.130 ;
        RECT  6.065 -0.130 6.615 0.325 ;
        RECT  0.385 -0.130 6.065 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 2.740 9.430 3.000 ;
        RECT  8.110 2.570 8.710 3.000 ;
        RECT  6.530 2.740 8.110 3.000 ;
        RECT  6.270 2.620 6.530 3.000 ;
        RECT  5.645 2.740 6.270 3.000 ;
        RECT  5.045 2.620 5.645 3.000 ;
        RECT  4.250 2.740 5.045 3.000 ;
        RECT  3.990 2.620 4.250 3.000 ;
        RECT  1.920 2.740 3.990 3.000 ;
        RECT  1.660 2.490 1.920 3.000 ;
        RECT  0.000 2.740 1.660 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.895 1.215 8.985 1.475 ;
        RECT  8.735 1.215 8.895 2.105 ;
        RECT  8.095 1.945 8.735 2.105 ;
        RECT  8.395 0.430 8.555 1.400 ;
        RECT  7.755 0.430 8.395 0.590 ;
        RECT  8.345 1.140 8.395 1.400 ;
        RECT  8.095 0.815 8.215 0.975 ;
        RECT  7.935 0.815 8.095 2.105 ;
        RECT  7.830 1.525 7.935 1.785 ;
        RECT  7.595 0.430 7.755 1.300 ;
        RECT  6.915 0.430 7.595 0.590 ;
        RECT  7.530 1.140 7.595 1.300 ;
        RECT  7.370 1.140 7.530 2.465 ;
        RECT  7.190 0.800 7.415 0.960 ;
        RECT  7.150 2.305 7.370 2.465 ;
        RECT  7.030 0.800 7.190 2.105 ;
        RECT  6.965 1.945 7.030 2.105 ;
        RECT  6.805 1.945 6.965 2.440 ;
        RECT  6.690 1.360 6.850 1.620 ;
        RECT  6.085 2.280 6.805 2.440 ;
        RECT  6.220 1.360 6.690 1.520 ;
        RECT  6.365 1.915 6.625 2.100 ;
        RECT  5.665 1.940 6.365 2.100 ;
        RECT  5.960 1.360 6.220 1.760 ;
        RECT  5.825 2.280 6.085 2.495 ;
        RECT  5.890 1.360 5.960 1.520 ;
        RECT  5.755 0.680 5.890 1.520 ;
        RECT  3.795 2.280 5.825 2.440 ;
        RECT  5.730 0.325 5.755 1.520 ;
        RECT  5.595 0.325 5.730 0.840 ;
        RECT  5.505 1.815 5.665 2.100 ;
        RECT  3.160 0.325 5.595 0.485 ;
        RECT  5.295 1.815 5.505 1.975 ;
        RECT  5.135 0.795 5.295 1.975 ;
        RECT  3.880 1.355 5.135 1.515 ;
        RECT  4.980 1.715 5.135 1.975 ;
        RECT  4.765 0.670 4.925 1.165 ;
        RECT  3.435 1.005 4.765 1.165 ;
        RECT  2.960 0.665 4.540 0.825 ;
        RECT  3.635 2.280 3.795 2.560 ;
        RECT  3.385 2.345 3.635 2.560 ;
        RECT  3.275 1.005 3.435 2.165 ;
        RECT  3.095 2.345 3.385 2.505 ;
        RECT  3.140 1.005 3.275 1.195 ;
        RECT  2.915 1.035 3.140 1.195 ;
        RECT  2.935 1.375 3.095 2.505 ;
        RECT  2.800 0.665 2.960 0.855 ;
        RECT  2.735 1.375 2.935 1.535 ;
        RECT  2.735 0.695 2.800 0.855 ;
        RECT  2.595 1.905 2.755 2.505 ;
        RECT  2.575 0.695 2.735 1.535 ;
        RECT  0.655 0.355 2.620 0.515 ;
        RECT  0.970 2.125 2.595 2.285 ;
        RECT  1.665 0.695 1.925 0.890 ;
        RECT  0.915 0.695 1.665 0.855 ;
        RECT  0.810 2.125 0.970 2.505 ;
        RECT  0.655 0.695 0.915 1.075 ;
        RECT  0.630 1.785 0.830 1.945 ;
        RECT  0.630 0.885 0.655 1.075 ;
        RECT  0.350 0.885 0.630 2.560 ;
    END
END SDFFQNX2MTH

MACRO SDFFQNX4MTH
    CLASS CORE ;
    FOREIGN SDFFQNX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.520 1.165 1.950 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.760 2.120 1.920 ;
        RECT  1.130 1.355 1.255 1.920 ;
        RECT  1.095 1.290 1.130 1.920 ;
        RECT  0.860 1.290 1.095 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.245 1.685 9.330 2.285 ;
        RECT  9.080 0.425 9.245 2.285 ;
        RECT  8.915 0.425 9.080 1.025 ;
        RECT  9.055 1.685 9.080 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.360 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.700 4.665 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.685 -0.130 9.840 0.130 ;
        RECT  9.425 -0.130 9.685 1.025 ;
        RECT  8.520 -0.130 9.425 0.130 ;
        RECT  7.920 -0.130 8.520 0.250 ;
        RECT  6.665 -0.130 7.920 0.130 ;
        RECT  6.065 -0.130 6.665 0.325 ;
        RECT  0.385 -0.130 6.065 0.130 ;
        RECT  0.125 -0.130 0.385 0.350 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 2.740 9.840 3.000 ;
        RECT  8.110 2.620 8.710 3.000 ;
        RECT  6.530 2.740 8.110 3.000 ;
        RECT  6.270 2.620 6.530 3.000 ;
        RECT  5.645 2.740 6.270 3.000 ;
        RECT  5.045 2.620 5.645 3.000 ;
        RECT  4.250 2.740 5.045 3.000 ;
        RECT  3.990 2.620 4.250 3.000 ;
        RECT  1.920 2.740 3.990 3.000 ;
        RECT  1.660 2.490 1.920 3.000 ;
        RECT  0.000 2.740 1.660 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.875 1.215 8.900 1.475 ;
        RECT  8.715 1.215 8.875 1.895 ;
        RECT  8.040 1.735 8.715 1.895 ;
        RECT  7.530 2.235 8.530 2.395 ;
        RECT  8.040 0.815 8.195 0.975 ;
        RECT  7.880 0.815 8.040 1.895 ;
        RECT  7.535 0.430 7.695 1.465 ;
        RECT  6.915 0.430 7.535 0.590 ;
        RECT  7.530 1.305 7.535 1.465 ;
        RECT  7.370 1.305 7.530 2.465 ;
        RECT  7.150 2.305 7.370 2.465 ;
        RECT  7.195 0.770 7.355 1.030 ;
        RECT  7.190 0.870 7.195 1.030 ;
        RECT  7.030 0.870 7.190 2.105 ;
        RECT  6.965 1.945 7.030 2.105 ;
        RECT  6.805 1.945 6.965 2.440 ;
        RECT  6.690 1.360 6.850 1.620 ;
        RECT  6.080 2.280 6.805 2.440 ;
        RECT  6.220 1.360 6.690 1.520 ;
        RECT  6.365 1.915 6.625 2.100 ;
        RECT  5.665 1.940 6.365 2.100 ;
        RECT  5.960 1.360 6.220 1.760 ;
        RECT  5.820 2.280 6.080 2.495 ;
        RECT  5.890 1.360 5.960 1.520 ;
        RECT  5.755 0.680 5.890 1.520 ;
        RECT  3.795 2.280 5.820 2.440 ;
        RECT  5.730 0.325 5.755 1.520 ;
        RECT  5.595 0.325 5.730 0.840 ;
        RECT  5.505 1.765 5.665 2.100 ;
        RECT  3.160 0.325 5.595 0.485 ;
        RECT  5.295 1.765 5.505 1.925 ;
        RECT  5.135 0.795 5.295 1.925 ;
        RECT  3.880 1.355 5.135 1.515 ;
        RECT  4.915 1.765 5.135 1.925 ;
        RECT  4.765 0.670 4.925 1.165 ;
        RECT  3.435 1.005 4.765 1.165 ;
        RECT  2.960 0.665 4.540 0.825 ;
        RECT  3.635 2.280 3.795 2.560 ;
        RECT  3.385 2.345 3.635 2.560 ;
        RECT  3.275 1.005 3.435 2.165 ;
        RECT  3.095 2.345 3.385 2.505 ;
        RECT  3.140 1.005 3.275 1.195 ;
        RECT  2.915 1.035 3.140 1.195 ;
        RECT  2.935 1.375 3.095 2.505 ;
        RECT  2.800 0.665 2.960 0.855 ;
        RECT  2.735 1.375 2.935 1.535 ;
        RECT  2.735 0.695 2.800 0.855 ;
        RECT  2.595 1.905 2.755 2.505 ;
        RECT  2.575 0.695 2.735 1.535 ;
        RECT  0.655 0.355 2.620 0.515 ;
        RECT  0.970 2.125 2.595 2.285 ;
        RECT  1.665 0.695 1.925 0.890 ;
        RECT  0.915 0.695 1.665 0.855 ;
        RECT  0.810 2.125 0.970 2.505 ;
        RECT  0.655 0.695 0.915 1.075 ;
        RECT  0.630 1.785 0.830 1.945 ;
        RECT  0.630 0.885 0.655 1.075 ;
        RECT  0.350 0.885 0.630 2.560 ;
    END
END SDFFQNX4MTH

MACRO SDFFQX1MTH
    CLASS CORE ;
    FOREIGN SDFFQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.435 1.160 1.950 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.760 2.155 1.920 ;
        RECT  1.130 1.355 1.255 1.920 ;
        RECT  1.095 1.290 1.130 1.920 ;
        RECT  0.915 1.290 1.095 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.300 1.290 9.330 1.580 ;
        RECT  9.040 0.705 9.300 2.015 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.360 1.580 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.700 4.665 1.990 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.010 -0.130 9.430 0.130 ;
        RECT  8.070 -0.130 9.010 0.250 ;
        RECT  6.710 -0.130 8.070 0.130 ;
        RECT  6.110 -0.130 6.710 0.350 ;
        RECT  0.405 -0.130 6.110 0.130 ;
        RECT  0.145 -0.130 0.405 0.300 ;
        RECT  0.000 -0.130 0.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.020 2.740 9.430 3.000 ;
        RECT  8.080 2.575 9.020 3.000 ;
        RECT  6.590 2.740 8.080 3.000 ;
        RECT  6.330 2.620 6.590 3.000 ;
        RECT  5.645 2.740 6.330 3.000 ;
        RECT  5.045 2.620 5.645 3.000 ;
        RECT  4.250 2.740 5.045 3.000 ;
        RECT  3.990 2.620 4.250 3.000 ;
        RECT  1.955 2.740 3.990 3.000 ;
        RECT  1.695 2.490 1.955 3.000 ;
        RECT  0.000 2.740 1.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.700 1.230 8.820 1.490 ;
        RECT  8.540 0.455 8.700 2.395 ;
        RECT  7.140 0.455 8.540 0.615 ;
        RECT  7.390 2.235 8.540 2.395 ;
        RECT  8.125 0.795 8.330 0.995 ;
        RECT  8.125 1.685 8.330 1.945 ;
        RECT  7.965 0.795 8.125 1.945 ;
        RECT  7.865 1.210 7.965 1.470 ;
        RECT  7.590 0.820 7.640 1.080 ;
        RECT  7.430 0.820 7.590 2.035 ;
        RECT  7.380 0.820 7.430 1.080 ;
        RECT  7.050 1.875 7.430 2.035 ;
        RECT  7.230 2.235 7.390 2.495 ;
        RECT  6.220 1.390 7.190 1.550 ;
        RECT  6.890 1.875 7.050 2.440 ;
        RECT  6.085 2.280 6.890 2.440 ;
        RECT  6.450 1.855 6.710 2.100 ;
        RECT  5.660 1.940 6.450 2.100 ;
        RECT  5.960 1.390 6.220 1.760 ;
        RECT  5.825 2.280 6.085 2.495 ;
        RECT  5.890 1.390 5.960 1.560 ;
        RECT  5.890 0.630 5.940 0.890 ;
        RECT  5.730 0.325 5.890 1.560 ;
        RECT  3.795 2.280 5.825 2.440 ;
        RECT  3.160 0.325 5.730 0.485 ;
        RECT  5.500 1.765 5.660 2.100 ;
        RECT  5.430 1.765 5.500 1.925 ;
        RECT  5.270 0.665 5.430 1.925 ;
        RECT  3.880 1.355 5.270 1.515 ;
        RECT  4.930 1.765 5.270 1.925 ;
        RECT  4.850 0.905 5.010 1.165 ;
        RECT  3.435 1.005 4.850 1.165 ;
        RECT  2.960 0.665 4.540 0.825 ;
        RECT  3.635 2.280 3.795 2.560 ;
        RECT  3.385 2.345 3.635 2.560 ;
        RECT  3.275 1.005 3.435 2.165 ;
        RECT  3.095 2.345 3.385 2.505 ;
        RECT  3.140 1.005 3.275 1.195 ;
        RECT  2.935 1.035 3.140 1.195 ;
        RECT  2.935 1.375 3.095 2.505 ;
        RECT  2.800 0.665 2.960 0.855 ;
        RECT  2.755 1.375 2.935 1.535 ;
        RECT  2.755 0.695 2.800 0.855 ;
        RECT  2.595 0.695 2.755 1.535 ;
        RECT  2.595 2.125 2.755 2.425 ;
        RECT  0.655 0.355 2.620 0.515 ;
        RECT  1.005 2.125 2.595 2.285 ;
        RECT  0.915 0.730 1.940 0.890 ;
        RECT  0.845 2.125 1.005 2.505 ;
        RECT  0.715 0.730 0.915 1.075 ;
        RECT  0.715 1.785 0.870 1.945 ;
        RECT  0.665 0.730 0.715 1.945 ;
        RECT  0.655 0.730 0.665 2.560 ;
        RECT  0.385 0.885 0.655 2.560 ;
    END
END SDFFQX1MTH

MACRO SDFFQX2MTH
    CLASS CORE ;
    FOREIGN SDFFQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.520 1.165 1.950 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.760 2.155 1.920 ;
        RECT  1.130 1.355 1.255 1.920 ;
        RECT  1.095 1.290 1.130 1.920 ;
        RECT  0.915 1.290 1.095 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.300 1.290 9.330 1.580 ;
        RECT  9.040 0.420 9.300 2.290 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.360 1.580 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.040 1.740 4.735 1.990 ;
        END
        AntennaGateArea 0.0871 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.670 -0.130 9.430 0.130 ;
        RECT  8.070 -0.130 8.670 0.250 ;
        RECT  6.475 -0.130 8.070 0.130 ;
        RECT  6.215 -0.130 6.475 0.350 ;
        RECT  0.385 -0.130 6.215 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.685 2.740 9.430 3.000 ;
        RECT  8.080 2.575 8.685 3.000 ;
        RECT  6.590 2.740 8.080 3.000 ;
        RECT  6.330 2.620 6.590 3.000 ;
        RECT  5.645 2.740 6.330 3.000 ;
        RECT  5.385 2.620 5.645 3.000 ;
        RECT  4.595 2.740 5.385 3.000 ;
        RECT  3.995 2.620 4.595 3.000 ;
        RECT  1.955 2.740 3.995 3.000 ;
        RECT  1.695 2.490 1.955 3.000 ;
        RECT  0.000 2.740 1.695 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.700 1.230 8.820 1.490 ;
        RECT  8.540 0.430 8.700 2.395 ;
        RECT  7.130 0.430 8.540 0.590 ;
        RECT  7.390 2.235 8.540 2.395 ;
        RECT  8.125 0.815 8.330 0.975 ;
        RECT  8.125 1.685 8.330 1.945 ;
        RECT  7.965 0.815 8.125 1.945 ;
        RECT  7.865 1.210 7.965 1.470 ;
        RECT  7.590 0.800 7.640 0.960 ;
        RECT  7.430 0.800 7.590 1.905 ;
        RECT  7.380 0.800 7.430 0.960 ;
        RECT  7.050 1.745 7.430 1.905 ;
        RECT  7.230 2.235 7.390 2.495 ;
        RECT  6.220 1.260 7.190 1.420 ;
        RECT  6.890 1.745 7.050 2.440 ;
        RECT  3.795 2.280 6.890 2.440 ;
        RECT  6.450 1.745 6.710 2.100 ;
        RECT  5.665 1.940 6.450 2.100 ;
        RECT  5.960 1.260 6.220 1.760 ;
        RECT  5.890 1.260 5.960 1.420 ;
        RECT  5.890 0.630 5.945 0.890 ;
        RECT  5.730 0.325 5.890 1.420 ;
        RECT  3.160 0.325 5.730 0.485 ;
        RECT  5.505 1.600 5.665 2.100 ;
        RECT  5.440 1.600 5.505 1.760 ;
        RECT  5.440 0.680 5.485 0.840 ;
        RECT  5.280 0.680 5.440 1.760 ;
        RECT  5.225 0.680 5.280 0.840 ;
        RECT  4.915 1.400 5.280 1.760 ;
        RECT  4.885 0.915 5.045 1.195 ;
        RECT  3.910 1.400 4.915 1.560 ;
        RECT  3.435 1.035 4.885 1.195 ;
        RECT  4.280 0.665 4.540 0.855 ;
        RECT  2.700 0.695 4.280 0.855 ;
        RECT  3.635 2.280 3.795 2.560 ;
        RECT  3.385 2.345 3.635 2.560 ;
        RECT  3.275 1.035 3.435 2.165 ;
        RECT  3.095 2.345 3.385 2.505 ;
        RECT  2.915 1.035 3.275 1.195 ;
        RECT  2.935 1.375 3.095 2.505 ;
        RECT  2.700 1.375 2.935 1.535 ;
        RECT  2.595 2.125 2.755 2.415 ;
        RECT  2.540 0.695 2.700 1.535 ;
        RECT  0.655 0.355 2.605 0.515 ;
        RECT  1.005 2.125 2.595 2.285 ;
        RECT  1.665 0.695 1.925 0.885 ;
        RECT  0.915 0.695 1.665 0.855 ;
        RECT  0.845 2.125 1.005 2.505 ;
        RECT  0.715 0.695 0.915 1.075 ;
        RECT  0.715 1.785 0.870 1.945 ;
        RECT  0.665 0.695 0.715 1.945 ;
        RECT  0.655 0.695 0.665 2.560 ;
        RECT  0.385 0.885 0.655 2.560 ;
    END
END SDFFQX2MTH

MACRO SDFFQX4MTH
    CLASS CORE ;
    FOREIGN SDFFQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.515 1.155 1.950 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.255 1.775 2.115 1.935 ;
        RECT  1.130 1.355 1.255 1.935 ;
        RECT  1.095 1.290 1.130 1.935 ;
        RECT  0.915 1.290 1.095 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.410 0.425 9.740 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 0.880 2.360 1.580 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.085 1.685 4.660 1.990 ;
        END
        AntennaGateArea 0.0988 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.130 -0.130 10.250 0.130 ;
        RECT  8.190 -0.130 9.130 0.295 ;
        RECT  6.360 -0.130 8.190 0.130 ;
        RECT  6.100 -0.130 6.360 0.300 ;
        RECT  0.390 -0.130 6.100 0.130 ;
        RECT  0.130 -0.130 0.390 0.300 ;
        RECT  0.000 -0.130 0.130 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.065 2.740 10.250 3.000 ;
        RECT  8.125 2.415 9.065 3.000 ;
        RECT  6.430 2.740 8.125 3.000 ;
        RECT  5.490 2.620 6.430 3.000 ;
        RECT  4.235 2.740 5.490 3.000 ;
        RECT  3.975 2.620 4.235 3.000 ;
        RECT  1.910 2.740 3.975 3.000 ;
        RECT  1.650 2.620 1.910 3.000 ;
        RECT  0.000 2.740 1.650 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.100 1.230 9.230 1.490 ;
        RECT  8.940 0.475 9.100 2.235 ;
        RECT  8.010 0.475 8.940 0.635 ;
        RECT  7.390 2.075 8.940 2.235 ;
        RECT  8.025 0.815 8.760 0.975 ;
        RECT  8.025 1.735 8.760 1.895 ;
        RECT  7.865 0.815 8.025 1.895 ;
        RECT  7.850 0.425 8.010 0.635 ;
        RECT  7.020 0.425 7.850 0.585 ;
        RECT  7.450 0.805 7.590 0.965 ;
        RECT  7.290 0.805 7.450 1.755 ;
        RECT  7.230 2.075 7.390 2.395 ;
        RECT  7.050 1.595 7.290 1.755 ;
        RECT  6.480 0.915 7.110 1.075 ;
        RECT  6.890 1.255 7.050 2.440 ;
        RECT  6.140 1.255 6.890 1.415 ;
        RECT  4.775 2.280 6.890 2.440 ;
        RECT  6.610 1.595 6.710 1.755 ;
        RECT  6.450 1.595 6.610 2.100 ;
        RECT  6.320 0.675 6.480 1.075 ;
        RECT  5.430 1.940 6.450 2.100 ;
        RECT  5.770 0.675 6.320 0.835 ;
        RECT  5.770 1.600 6.220 1.760 ;
        RECT  5.980 1.065 6.140 1.415 ;
        RECT  5.610 0.325 5.770 1.760 ;
        RECT  3.160 0.325 5.610 0.485 ;
        RECT  5.270 0.665 5.430 2.100 ;
        RECT  5.090 1.345 5.270 2.100 ;
        RECT  3.865 1.345 5.090 1.505 ;
        RECT  4.965 1.755 5.090 2.100 ;
        RECT  4.890 0.905 5.060 1.165 ;
        RECT  3.395 1.005 4.890 1.165 ;
        RECT  4.515 2.280 4.775 2.465 ;
        RECT  2.945 0.665 4.540 0.825 ;
        RECT  3.795 2.280 4.515 2.440 ;
        RECT  3.635 2.280 3.795 2.545 ;
        RECT  3.385 2.345 3.635 2.545 ;
        RECT  3.235 1.005 3.395 2.165 ;
        RECT  3.055 2.345 3.385 2.505 ;
        RECT  3.140 1.005 3.235 1.195 ;
        RECT  2.915 1.035 3.140 1.195 ;
        RECT  2.895 1.375 3.055 2.505 ;
        RECT  2.785 0.665 2.945 0.855 ;
        RECT  2.700 1.375 2.895 1.535 ;
        RECT  2.700 0.695 2.785 0.855 ;
        RECT  2.555 2.240 2.715 2.505 ;
        RECT  2.540 0.695 2.700 1.535 ;
        RECT  0.655 0.355 2.605 0.515 ;
        RECT  0.960 2.240 2.555 2.400 ;
        RECT  1.665 0.695 1.925 0.885 ;
        RECT  0.915 0.695 1.665 0.855 ;
        RECT  0.800 2.240 0.960 2.505 ;
        RECT  0.655 0.695 0.915 1.075 ;
        RECT  0.620 1.785 0.820 1.945 ;
        RECT  0.590 0.915 0.655 1.075 ;
        RECT  0.590 1.785 0.620 2.560 ;
        RECT  0.360 0.915 0.590 2.560 ;
    END
END SDFFQX4MTH

MACRO SDFFRHQX1MTH
    CLASS CORE ;
    FOREIGN SDFFRHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 1.280 5.270 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.170 0.800 5.330 1.100 ;
        RECT  4.435 0.880 5.170 1.040 ;
        RECT  3.930 0.880 4.435 1.170 ;
        RECT  3.670 0.880 3.930 1.200 ;
        END
        AntennaGateArea 0.1118 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.350 1.025 10.610 1.635 ;
        END
        AntennaGateArea 0.143 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.580 1.290 12.610 1.580 ;
        RECT  12.400 0.725 12.580 2.070 ;
        RECT  12.375 0.725 12.400 0.985 ;
        RECT  12.375 1.765 12.400 2.025 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.510 0.880 2.770 1.330 ;
        RECT  2.150 0.880 2.510 1.180 ;
        END
        AntennaGateArea 0.1105 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.105 0.760 1.660 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.560 -0.130 12.710 0.130 ;
        RECT  12.300 -0.130 12.560 0.300 ;
        RECT  12.045 -0.130 12.300 0.130 ;
        RECT  11.785 -0.130 12.045 0.490 ;
        RECT  11.375 -0.130 11.785 0.130 ;
        RECT  10.775 -0.130 11.375 0.485 ;
        RECT  8.375 -0.130 10.775 0.130 ;
        RECT  7.775 -0.130 8.375 0.450 ;
        RECT  4.650 -0.130 7.775 0.130 ;
        RECT  4.390 -0.130 4.650 0.250 ;
        RECT  2.485 -0.130 4.390 0.130 ;
        RECT  2.285 -0.130 2.485 0.700 ;
        RECT  0.635 -0.130 2.285 0.130 ;
        RECT  0.375 -0.130 0.635 0.300 ;
        RECT  0.000 -0.130 0.375 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.890 2.740 12.710 3.000 ;
        RECT  11.630 2.415 11.890 3.000 ;
        RECT  10.145 2.740 11.630 3.000 ;
        RECT  9.885 2.295 10.145 3.000 ;
        RECT  8.650 2.740 9.885 3.000 ;
        RECT  8.390 2.620 8.650 3.000 ;
        RECT  7.655 2.740 8.390 3.000 ;
        RECT  7.395 2.620 7.655 3.000 ;
        RECT  1.960 2.740 7.395 3.000 ;
        RECT  1.700 2.570 1.960 3.000 ;
        RECT  0.815 2.740 1.700 3.000 ;
        RECT  0.215 2.455 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.025 1.230 12.220 1.490 ;
        RECT  11.865 1.230 12.025 2.235 ;
        RECT  11.720 1.230 11.865 1.490 ;
        RECT  11.450 2.075 11.865 2.235 ;
        RECT  11.515 1.735 11.615 1.895 ;
        RECT  11.355 0.740 11.515 1.895 ;
        RECT  11.290 2.075 11.450 2.455 ;
        RECT  11.310 0.740 11.355 1.455 ;
        RECT  11.145 1.195 11.310 1.455 ;
        RECT  10.495 2.295 11.290 2.455 ;
        RECT  10.790 0.685 10.950 2.115 ;
        RECT  10.555 0.685 10.790 0.845 ;
        RECT  10.715 1.855 10.790 2.115 ;
        RECT  10.395 0.310 10.555 0.845 ;
        RECT  10.335 1.955 10.495 2.455 ;
        RECT  8.790 0.310 10.395 0.470 ;
        RECT  10.170 1.955 10.335 2.115 ;
        RECT  10.010 0.800 10.170 2.115 ;
        RECT  9.835 0.800 10.010 0.960 ;
        RECT  9.935 1.735 10.010 2.115 ;
        RECT  9.575 0.700 9.835 0.960 ;
        RECT  9.705 1.250 9.830 1.530 ;
        RECT  9.670 1.250 9.705 2.440 ;
        RECT  9.545 1.370 9.670 2.440 ;
        RECT  7.060 2.280 9.545 2.440 ;
        RECT  9.205 0.690 9.365 2.000 ;
        RECT  8.970 0.690 9.205 0.850 ;
        RECT  9.185 1.840 9.205 2.000 ;
        RECT  9.025 1.840 9.185 2.100 ;
        RECT  7.430 1.940 9.025 2.100 ;
        RECT  8.235 1.075 9.010 1.335 ;
        RECT  8.630 0.310 8.790 0.810 ;
        RECT  7.380 0.650 8.630 0.810 ;
        RECT  7.975 0.990 8.235 1.755 ;
        RECT  6.720 0.990 7.975 1.150 ;
        RECT  7.270 1.400 7.430 2.100 ;
        RECT  7.220 0.365 7.380 0.810 ;
        RECT  6.040 0.650 7.220 0.810 ;
        RECT  6.900 2.280 7.060 2.560 ;
        RECT  4.990 0.310 6.915 0.470 ;
        RECT  6.380 2.400 6.900 2.560 ;
        RECT  6.560 0.990 6.720 2.210 ;
        RECT  6.220 1.065 6.380 2.560 ;
        RECT  2.335 2.400 6.220 2.560 ;
        RECT  5.880 0.650 6.040 2.220 ;
        RECT  2.675 2.060 5.880 2.220 ;
        RECT  5.540 0.650 5.700 1.880 ;
        RECT  4.545 1.720 5.540 1.880 ;
        RECT  4.830 0.310 4.990 0.695 ;
        RECT  3.490 0.535 4.830 0.695 ;
        RECT  4.385 1.350 4.545 1.880 ;
        RECT  4.175 1.350 4.385 1.510 ;
        RECT  3.980 1.720 4.205 1.880 ;
        RECT  3.820 1.380 3.980 1.880 ;
        RECT  3.490 1.380 3.820 1.540 ;
        RECT  3.145 1.720 3.635 1.880 ;
        RECT  3.330 0.535 3.490 1.540 ;
        RECT  2.985 0.530 3.145 1.880 ;
        RECT  2.805 0.530 2.985 0.690 ;
        RECT  2.855 1.550 2.985 1.880 ;
        RECT  2.515 1.600 2.675 2.220 ;
        RECT  1.925 1.600 2.515 1.760 ;
        RECT  2.175 2.110 2.335 2.560 ;
        RECT  1.105 2.110 2.175 2.270 ;
        RECT  0.975 0.310 2.105 0.470 ;
        RECT  1.765 0.680 1.925 1.760 ;
        RECT  1.665 0.680 1.765 0.840 ;
        RECT  1.445 1.600 1.765 1.760 ;
        RECT  1.285 1.470 1.445 1.760 ;
        RECT  1.315 0.680 1.415 0.840 ;
        RECT  1.155 0.680 1.315 1.280 ;
        RECT  1.105 1.120 1.155 1.280 ;
        RECT  0.945 1.120 1.105 2.270 ;
        RECT  0.815 0.310 0.975 0.925 ;
        RECT  0.360 0.765 0.815 0.925 ;
        RECT  0.330 0.665 0.360 0.925 ;
        RECT  0.330 1.860 0.360 2.120 ;
        RECT  0.170 0.665 0.330 2.120 ;
    END
END SDFFRHQX1MTH

MACRO SDFFRHQX2MTH
    CLASS CORE ;
    FOREIGN SDFFRHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.730 1.280 5.325 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.170 0.840 5.330 1.100 ;
        RECT  4.410 0.880 5.170 1.040 ;
        RECT  3.930 0.880 4.410 1.170 ;
        RECT  3.670 0.880 3.930 1.200 ;
        END
        AntennaGateArea 0.1274 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.120 1.025 11.380 1.680 ;
        RECT  11.080 1.420 11.120 1.680 ;
        END
        AntennaGateArea 0.1664 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.190 0.385 13.430 2.405 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 0.880 2.780 1.180 ;
        RECT  2.560 0.880 2.720 1.380 ;
        RECT  2.150 0.880 2.560 1.180 ;
        END
        AntennaGateArea 0.0923 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.105 0.760 1.660 ;
        END
        AntennaGateArea 0.143 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.895 -0.130 13.530 0.130 ;
        RECT  12.635 -0.130 12.895 0.985 ;
        RECT  12.055 -0.130 12.635 0.130 ;
        RECT  11.455 -0.130 12.055 0.480 ;
        RECT  8.680 -0.130 11.455 0.130 ;
        RECT  7.740 -0.130 8.680 0.460 ;
        RECT  4.650 -0.130 7.740 0.130 ;
        RECT  4.390 -0.130 4.650 0.250 ;
        RECT  2.485 -0.130 4.390 0.130 ;
        RECT  2.285 -0.130 2.485 0.700 ;
        RECT  0.685 -0.130 2.285 0.130 ;
        RECT  0.185 -0.130 0.685 0.300 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.845 2.740 13.530 3.000 ;
        RECT  12.245 2.415 12.845 3.000 ;
        RECT  10.930 2.740 12.245 3.000 ;
        RECT  10.670 2.295 10.930 3.000 ;
        RECT  8.955 2.740 10.670 3.000 ;
        RECT  8.695 2.620 8.955 3.000 ;
        RECT  7.855 2.740 8.695 3.000 ;
        RECT  7.595 2.620 7.855 3.000 ;
        RECT  1.790 2.740 7.595 3.000 ;
        RECT  1.630 2.570 1.790 3.000 ;
        RECT  0.815 2.740 1.630 3.000 ;
        RECT  0.215 2.350 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.745 1.230 13.010 1.490 ;
        RECT  12.585 1.230 12.745 2.235 ;
        RECT  12.450 1.230 12.585 1.490 ;
        RECT  12.065 2.075 12.585 2.235 ;
        RECT  12.250 1.735 12.405 1.895 ;
        RECT  12.090 0.765 12.250 1.895 ;
        RECT  12.070 0.765 12.090 1.395 ;
        RECT  11.900 1.135 12.070 1.395 ;
        RECT  11.905 2.075 12.065 2.455 ;
        RECT  11.280 2.295 11.905 2.455 ;
        RECT  11.560 0.685 11.720 2.115 ;
        RECT  11.275 0.685 11.560 0.845 ;
        RECT  11.505 1.855 11.560 2.115 ;
        RECT  11.120 1.955 11.280 2.455 ;
        RECT  11.115 0.310 11.275 0.845 ;
        RECT  10.900 1.955 11.120 2.115 ;
        RECT  10.075 0.310 11.115 0.470 ;
        RECT  10.740 0.650 10.900 2.115 ;
        RECT  10.255 0.650 10.740 0.810 ;
        RECT  10.070 1.955 10.740 2.115 ;
        RECT  10.300 1.470 10.560 1.775 ;
        RECT  9.735 1.470 10.300 1.630 ;
        RECT  9.915 0.310 10.075 1.145 ;
        RECT  9.910 1.815 10.070 2.115 ;
        RECT  9.115 0.310 9.915 0.470 ;
        RECT  9.760 1.815 9.910 1.975 ;
        RECT  9.480 2.185 9.740 2.440 ;
        RECT  9.580 0.650 9.735 1.630 ;
        RECT  9.575 0.650 9.580 1.980 ;
        RECT  9.405 0.650 9.575 0.810 ;
        RECT  9.420 1.470 9.575 1.980 ;
        RECT  7.410 2.280 9.480 2.440 ;
        RECT  9.300 1.720 9.420 1.980 ;
        RECT  9.155 0.990 9.315 1.315 ;
        RECT  9.140 1.720 9.300 2.100 ;
        RECT  8.405 0.990 9.155 1.150 ;
        RECT  7.705 1.940 9.140 2.100 ;
        RECT  8.955 0.310 9.115 0.810 ;
        RECT  7.380 0.650 8.955 0.810 ;
        RECT  8.405 1.480 8.575 1.710 ;
        RECT  8.145 0.990 8.405 1.710 ;
        RECT  7.065 0.990 8.145 1.150 ;
        RECT  7.975 1.480 8.145 1.710 ;
        RECT  7.545 1.455 7.705 2.100 ;
        RECT  7.250 2.280 7.410 2.560 ;
        RECT  7.220 0.365 7.380 0.810 ;
        RECT  6.715 2.400 7.250 2.560 ;
        RECT  6.040 0.650 7.220 0.810 ;
        RECT  6.905 0.990 7.065 2.210 ;
        RECT  4.990 0.310 6.915 0.470 ;
        RECT  6.555 1.165 6.715 2.560 ;
        RECT  6.380 1.165 6.555 1.325 ;
        RECT  2.335 2.400 6.555 2.560 ;
        RECT  6.220 1.065 6.380 1.325 ;
        RECT  6.040 1.545 6.355 1.805 ;
        RECT  5.880 0.650 6.040 2.220 ;
        RECT  2.675 2.060 5.880 2.220 ;
        RECT  5.540 0.650 5.700 1.880 ;
        RECT  4.545 1.720 5.540 1.880 ;
        RECT  4.830 0.310 4.990 0.695 ;
        RECT  3.490 0.535 4.830 0.695 ;
        RECT  4.385 1.350 4.545 1.880 ;
        RECT  4.160 1.350 4.385 1.510 ;
        RECT  3.980 1.720 4.205 1.880 ;
        RECT  3.820 1.380 3.980 1.880 ;
        RECT  3.490 1.380 3.820 1.540 ;
        RECT  3.145 1.720 3.635 1.880 ;
        RECT  3.330 0.535 3.490 1.540 ;
        RECT  2.985 0.530 3.145 1.880 ;
        RECT  2.805 0.530 2.985 0.690 ;
        RECT  2.855 1.620 2.985 1.880 ;
        RECT  2.515 1.585 2.675 2.220 ;
        RECT  2.095 1.585 2.515 1.745 ;
        RECT  2.175 2.055 2.335 2.560 ;
        RECT  1.665 2.055 2.175 2.215 ;
        RECT  1.025 0.310 2.105 0.470 ;
        RECT  1.925 1.585 2.095 1.845 ;
        RECT  1.835 0.700 1.925 1.845 ;
        RECT  1.765 0.700 1.835 1.745 ;
        RECT  1.665 0.700 1.765 0.860 ;
        RECT  1.445 1.585 1.765 1.745 ;
        RECT  1.405 2.055 1.665 2.270 ;
        RECT  1.285 1.470 1.445 1.745 ;
        RECT  1.105 2.055 1.405 2.215 ;
        RECT  1.205 0.665 1.365 1.280 ;
        RECT  1.105 1.120 1.205 1.280 ;
        RECT  0.945 1.120 1.105 2.215 ;
        RECT  0.865 0.310 1.025 0.925 ;
        RECT  0.370 0.765 0.865 0.925 ;
        RECT  0.330 0.665 0.370 0.925 ;
        RECT  0.330 1.840 0.370 2.100 ;
        RECT  0.170 0.665 0.330 2.100 ;
    END
END SDFFRHQX2MTH

MACRO SDFFRHQX4MTH
    CLASS CORE ;
    FOREIGN SDFFRHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.940 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 1.330 5.280 1.540 ;
        RECT  4.735 1.015 4.945 1.540 ;
        RECT  4.635 1.015 4.735 1.175 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.170 0.675 5.330 1.150 ;
        RECT  4.410 0.675 5.170 0.835 ;
        RECT  4.200 0.675 4.410 1.170 ;
        RECT  3.930 1.010 4.200 1.170 ;
        RECT  3.670 1.010 3.930 1.200 ;
        END
        AntennaGateArea 0.1274 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.120 1.085 11.380 1.635 ;
        RECT  11.080 1.375 11.120 1.635 ;
        END
        AntennaGateArea 0.1703 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.400 1.700 13.430 1.990 ;
        RECT  13.160 0.385 13.400 2.405 ;
        RECT  13.095 0.385 13.160 0.985 ;
        RECT  13.125 1.805 13.160 2.405 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 0.880 2.780 1.180 ;
        RECT  2.560 0.880 2.720 1.380 ;
        RECT  2.150 0.880 2.560 1.180 ;
        END
        AntennaGateArea 0.1664 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.105 0.760 1.660 ;
        END
        AntennaGateArea 0.1612 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.765 -0.130 13.940 0.130 ;
        RECT  13.605 -0.130 13.765 0.985 ;
        RECT  12.765 -0.130 13.605 0.130 ;
        RECT  12.505 -0.130 12.765 0.515 ;
        RECT  12.020 -0.130 12.505 0.130 ;
        RECT  11.420 -0.130 12.020 0.515 ;
        RECT  8.685 -0.130 11.420 0.130 ;
        RECT  7.745 -0.130 8.685 0.460 ;
        RECT  3.645 -0.130 7.745 0.130 ;
        RECT  3.485 -0.130 3.645 0.300 ;
        RECT  2.485 -0.130 3.485 0.130 ;
        RECT  2.285 -0.130 2.485 0.680 ;
        RECT  0.685 -0.130 2.285 0.130 ;
        RECT  0.185 -0.130 0.685 0.300 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.745 2.740 13.940 3.000 ;
        RECT  12.245 2.415 12.745 3.000 ;
        RECT  10.930 2.740 12.245 3.000 ;
        RECT  10.670 2.295 10.930 3.000 ;
        RECT  8.955 2.740 10.670 3.000 ;
        RECT  8.695 2.620 8.955 3.000 ;
        RECT  7.855 2.740 8.695 3.000 ;
        RECT  7.595 2.620 7.855 3.000 ;
        RECT  1.960 2.740 7.595 3.000 ;
        RECT  1.800 2.570 1.960 3.000 ;
        RECT  0.835 2.740 1.800 3.000 ;
        RECT  0.235 2.390 0.835 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.745 1.230 12.980 1.490 ;
        RECT  12.585 1.230 12.745 2.235 ;
        RECT  12.480 1.230 12.585 1.490 ;
        RECT  12.065 2.075 12.585 2.235 ;
        RECT  12.250 1.735 12.360 1.895 ;
        RECT  12.090 0.765 12.250 1.895 ;
        RECT  12.070 0.765 12.090 1.395 ;
        RECT  11.900 1.135 12.070 1.395 ;
        RECT  11.905 2.075 12.065 2.455 ;
        RECT  11.270 2.295 11.905 2.455 ;
        RECT  11.560 0.745 11.720 2.115 ;
        RECT  11.240 0.745 11.560 0.905 ;
        RECT  11.460 1.855 11.560 2.115 ;
        RECT  11.110 1.955 11.270 2.455 ;
        RECT  11.080 0.310 11.240 0.905 ;
        RECT  10.900 1.955 11.110 2.115 ;
        RECT  9.995 0.310 11.080 0.470 ;
        RECT  10.740 0.650 10.900 2.115 ;
        RECT  10.175 0.650 10.740 0.810 ;
        RECT  10.070 1.955 10.740 2.115 ;
        RECT  10.300 1.470 10.560 1.775 ;
        RECT  9.655 1.470 10.300 1.630 ;
        RECT  9.910 1.815 10.070 2.115 ;
        RECT  9.835 0.310 9.995 1.145 ;
        RECT  9.760 1.815 9.910 1.975 ;
        RECT  9.095 0.310 9.835 0.470 ;
        RECT  9.480 2.185 9.740 2.440 ;
        RECT  9.580 0.650 9.655 1.630 ;
        RECT  9.495 0.650 9.580 1.980 ;
        RECT  9.275 0.650 9.495 0.810 ;
        RECT  9.420 1.470 9.495 1.980 ;
        RECT  7.415 2.280 9.480 2.440 ;
        RECT  9.300 1.720 9.420 1.980 ;
        RECT  9.155 0.990 9.315 1.315 ;
        RECT  9.140 1.720 9.300 2.100 ;
        RECT  8.575 0.990 9.155 1.150 ;
        RECT  7.705 1.940 9.140 2.100 ;
        RECT  8.935 0.310 9.095 0.810 ;
        RECT  7.380 0.650 8.935 0.810 ;
        RECT  7.975 0.990 8.575 1.545 ;
        RECT  7.065 0.990 7.975 1.150 ;
        RECT  7.545 1.400 7.705 2.100 ;
        RECT  7.255 2.280 7.415 2.560 ;
        RECT  7.220 0.365 7.380 0.810 ;
        RECT  6.715 2.400 7.255 2.560 ;
        RECT  6.040 0.650 7.220 0.810 ;
        RECT  6.905 0.990 7.065 2.210 ;
        RECT  3.985 0.310 6.915 0.470 ;
        RECT  6.555 1.165 6.715 2.560 ;
        RECT  6.380 1.165 6.555 1.325 ;
        RECT  2.300 2.400 6.555 2.560 ;
        RECT  6.220 1.065 6.380 1.325 ;
        RECT  6.040 1.545 6.355 1.805 ;
        RECT  5.880 0.650 6.040 2.220 ;
        RECT  2.670 2.060 5.880 2.220 ;
        RECT  5.540 0.650 5.700 1.880 ;
        RECT  4.515 1.720 5.540 1.880 ;
        RECT  4.355 1.350 4.515 1.880 ;
        RECT  4.155 1.350 4.355 1.510 ;
        RECT  3.975 1.720 4.175 1.880 ;
        RECT  3.825 0.310 3.985 0.800 ;
        RECT  3.815 1.380 3.975 1.880 ;
        RECT  3.490 0.640 3.825 0.800 ;
        RECT  3.490 1.380 3.815 1.540 ;
        RECT  3.145 1.720 3.635 1.880 ;
        RECT  3.330 0.640 3.490 1.540 ;
        RECT  2.985 0.530 3.145 1.880 ;
        RECT  2.775 0.530 2.985 0.690 ;
        RECT  2.855 1.620 2.985 1.880 ;
        RECT  2.510 1.630 2.670 2.220 ;
        RECT  1.960 1.630 2.510 1.790 ;
        RECT  2.140 2.055 2.300 2.560 ;
        RECT  1.685 2.055 2.140 2.215 ;
        RECT  1.025 0.310 2.105 0.470 ;
        RECT  1.800 0.700 1.960 1.790 ;
        RECT  1.665 0.700 1.800 0.860 ;
        RECT  1.465 1.630 1.800 1.790 ;
        RECT  1.425 2.055 1.685 2.270 ;
        RECT  1.305 1.470 1.465 1.790 ;
        RECT  1.105 2.055 1.425 2.215 ;
        RECT  1.205 0.660 1.365 1.280 ;
        RECT  1.105 1.120 1.205 1.280 ;
        RECT  0.945 1.120 1.105 2.215 ;
        RECT  0.865 0.310 1.025 0.820 ;
        RECT  0.375 0.660 0.865 0.820 ;
        RECT  0.330 0.660 0.375 0.920 ;
        RECT  0.330 1.840 0.375 2.100 ;
        RECT  0.170 0.660 0.330 2.100 ;
    END
END SDFFRHQX4MTH

MACRO SDFFRHQX8MTH
    CLASS CORE ;
    FOREIGN SDFFRHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.760 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 1.330 5.280 1.540 ;
        RECT  4.735 1.015 4.945 1.540 ;
        RECT  4.635 1.015 4.735 1.175 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.170 0.675 5.330 1.150 ;
        RECT  4.410 0.675 5.170 0.835 ;
        RECT  4.200 0.675 4.410 1.170 ;
        RECT  3.930 1.010 4.200 1.170 ;
        RECT  3.670 1.010 3.930 1.200 ;
        END
        AntennaGateArea 0.1274 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.120 1.085 11.380 1.635 ;
        RECT  11.080 1.375 11.120 1.635 ;
        END
        AntennaGateArea 0.1703 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.125 1.085 14.165 2.405 ;
        RECT  13.815 0.385 14.125 2.405 ;
        RECT  13.775 0.385 13.815 1.785 ;
        RECT  13.410 1.085 13.775 1.785 ;
        RECT  13.060 0.385 13.410 2.405 ;
        RECT  12.930 0.385 13.060 0.985 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.720 0.880 2.780 1.180 ;
        RECT  2.560 0.880 2.720 1.380 ;
        RECT  2.150 0.880 2.560 1.180 ;
        END
        AntennaGateArea 0.1664 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.105 0.760 1.660 ;
        END
        AntennaGateArea 0.1612 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.635 -0.130 14.760 0.130 ;
        RECT  14.375 -0.130 14.635 0.985 ;
        RECT  12.645 -0.130 14.375 0.130 ;
        RECT  12.385 -0.130 12.645 0.515 ;
        RECT  12.130 -0.130 12.385 0.130 ;
        RECT  11.530 -0.130 12.130 0.515 ;
        RECT  8.685 -0.130 11.530 0.130 ;
        RECT  7.745 -0.130 8.685 0.460 ;
        RECT  3.645 -0.130 7.745 0.130 ;
        RECT  3.485 -0.130 3.645 0.300 ;
        RECT  2.485 -0.130 3.485 0.130 ;
        RECT  2.285 -0.130 2.485 0.680 ;
        RECT  0.685 -0.130 2.285 0.130 ;
        RECT  0.185 -0.130 0.685 0.300 ;
        RECT  0.000 -0.130 0.185 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.660 2.740 14.760 3.000 ;
        RECT  12.240 2.415 12.660 3.000 ;
        RECT  10.885 2.740 12.240 3.000 ;
        RECT  10.625 2.295 10.885 3.000 ;
        RECT  8.955 2.740 10.625 3.000 ;
        RECT  8.695 2.620 8.955 3.000 ;
        RECT  7.855 2.740 8.695 3.000 ;
        RECT  7.595 2.620 7.855 3.000 ;
        RECT  1.960 2.740 7.595 3.000 ;
        RECT  1.800 2.570 1.960 3.000 ;
        RECT  0.835 2.740 1.800 3.000 ;
        RECT  0.235 2.390 0.835 3.000 ;
        RECT  0.000 2.740 0.235 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.700 1.230 12.880 1.490 ;
        RECT  12.540 1.230 12.700 2.235 ;
        RECT  12.380 1.230 12.540 1.490 ;
        RECT  12.060 2.075 12.540 2.235 ;
        RECT  12.115 1.735 12.315 1.895 ;
        RECT  12.115 0.765 12.170 1.025 ;
        RECT  11.955 0.765 12.115 1.895 ;
        RECT  11.900 2.075 12.060 2.455 ;
        RECT  11.900 1.135 11.955 1.395 ;
        RECT  11.235 2.295 11.900 2.455 ;
        RECT  11.560 0.745 11.720 2.115 ;
        RECT  11.245 0.745 11.560 0.905 ;
        RECT  11.415 1.855 11.560 2.115 ;
        RECT  11.085 0.310 11.245 0.905 ;
        RECT  11.075 1.955 11.235 2.455 ;
        RECT  10.045 0.310 11.085 0.470 ;
        RECT  10.855 1.955 11.075 2.115 ;
        RECT  10.695 0.650 10.855 2.115 ;
        RECT  10.225 0.650 10.695 0.810 ;
        RECT  10.070 1.955 10.695 2.115 ;
        RECT  10.255 1.470 10.515 1.775 ;
        RECT  9.705 1.470 10.255 1.630 ;
        RECT  9.910 1.815 10.070 2.115 ;
        RECT  9.885 0.310 10.045 1.145 ;
        RECT  9.715 1.815 9.910 1.975 ;
        RECT  9.095 0.310 9.885 0.470 ;
        RECT  9.545 0.650 9.705 1.630 ;
        RECT  9.375 2.185 9.635 2.440 ;
        RECT  9.275 0.650 9.545 0.810 ;
        RECT  9.535 1.470 9.545 1.630 ;
        RECT  9.375 1.470 9.535 1.980 ;
        RECT  9.195 1.720 9.375 1.980 ;
        RECT  7.415 2.280 9.375 2.440 ;
        RECT  9.155 0.990 9.315 1.290 ;
        RECT  9.035 1.720 9.195 2.100 ;
        RECT  8.575 0.990 9.155 1.150 ;
        RECT  8.935 0.310 9.095 0.810 ;
        RECT  7.705 1.940 9.035 2.100 ;
        RECT  7.380 0.650 8.935 0.810 ;
        RECT  7.975 0.990 8.575 1.545 ;
        RECT  7.065 0.990 7.975 1.150 ;
        RECT  7.545 1.400 7.705 2.100 ;
        RECT  7.255 2.280 7.415 2.560 ;
        RECT  7.220 0.365 7.380 0.810 ;
        RECT  6.715 2.400 7.255 2.560 ;
        RECT  6.040 0.650 7.220 0.810 ;
        RECT  6.905 0.990 7.065 2.210 ;
        RECT  3.985 0.310 6.915 0.470 ;
        RECT  6.555 1.165 6.715 2.560 ;
        RECT  6.380 1.165 6.555 1.325 ;
        RECT  2.300 2.400 6.555 2.560 ;
        RECT  6.220 1.065 6.380 1.325 ;
        RECT  6.040 1.545 6.355 1.805 ;
        RECT  5.880 0.650 6.040 2.220 ;
        RECT  2.670 2.060 5.880 2.220 ;
        RECT  5.540 0.650 5.700 1.880 ;
        RECT  4.515 1.720 5.540 1.880 ;
        RECT  4.355 1.350 4.515 1.880 ;
        RECT  4.155 1.350 4.355 1.510 ;
        RECT  3.975 1.720 4.175 1.880 ;
        RECT  3.825 0.310 3.985 0.800 ;
        RECT  3.815 1.380 3.975 1.880 ;
        RECT  3.490 0.640 3.825 0.800 ;
        RECT  3.490 1.380 3.815 1.540 ;
        RECT  3.145 1.720 3.635 1.880 ;
        RECT  3.330 0.640 3.490 1.540 ;
        RECT  2.985 0.530 3.145 1.880 ;
        RECT  2.775 0.530 2.985 0.690 ;
        RECT  2.855 1.620 2.985 1.880 ;
        RECT  2.510 1.630 2.670 2.220 ;
        RECT  1.960 1.630 2.510 1.790 ;
        RECT  2.140 2.055 2.300 2.560 ;
        RECT  1.685 2.055 2.140 2.215 ;
        RECT  1.025 0.310 2.105 0.470 ;
        RECT  1.800 0.700 1.960 1.790 ;
        RECT  1.665 0.700 1.800 0.860 ;
        RECT  1.465 1.630 1.800 1.790 ;
        RECT  1.425 2.055 1.685 2.270 ;
        RECT  1.305 1.470 1.465 1.790 ;
        RECT  1.105 2.055 1.425 2.215 ;
        RECT  1.205 0.660 1.365 1.280 ;
        RECT  1.105 1.120 1.205 1.280 ;
        RECT  0.945 1.120 1.105 2.215 ;
        RECT  0.865 0.310 1.025 0.820 ;
        RECT  0.375 0.660 0.865 0.820 ;
        RECT  0.330 0.660 0.375 0.920 ;
        RECT  0.330 1.840 0.375 2.100 ;
        RECT  0.170 0.660 0.330 2.100 ;
    END
END SDFFRHQX8MTH

MACRO SDFFRQX1MTH
    CLASS CORE ;
    FOREIGN SDFFRQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.120 2.770 1.785 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 1.465 1.610 1.725 ;
        RECT  0.760 1.465 1.350 1.630 ;
        RECT  0.465 1.275 0.760 1.630 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.190 1.040 9.735 1.200 ;
        RECT  9.030 0.325 9.190 1.200 ;
        RECT  7.765 0.325 9.030 0.485 ;
        RECT  7.605 0.325 7.765 1.145 ;
        RECT  7.165 0.920 7.605 1.145 ;
        RECT  6.895 0.920 7.165 1.115 ;
        RECT  6.735 0.310 6.895 1.115 ;
        RECT  3.745 0.310 6.735 0.470 ;
        RECT  3.585 0.310 3.745 0.645 ;
        RECT  3.295 0.485 3.585 0.645 ;
        RECT  3.230 0.485 3.295 1.380 ;
        RECT  3.135 0.485 3.230 1.785 ;
        RECT  3.070 1.185 3.135 1.785 ;
        END
        AntennaGateArea 0.1586 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.170 0.705 11.380 2.015 ;
        RECT  11.095 0.705 11.170 0.995 ;
        RECT  11.095 1.755 11.170 2.015 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 2.150 1.220 2.545 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 1.330 4.450 1.540 ;
        RECT  3.830 1.220 3.990 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 -0.130 11.480 0.130 ;
        RECT  10.345 -0.130 10.945 0.300 ;
        RECT  9.970 -0.130 10.345 0.130 ;
        RECT  9.370 -0.130 9.970 0.300 ;
        RECT  7.425 -0.130 9.370 0.130 ;
        RECT  7.195 -0.130 7.425 0.740 ;
        RECT  3.405 -0.130 7.195 0.130 ;
        RECT  2.905 -0.130 3.405 0.300 ;
        RECT  0.725 -0.130 2.905 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.730 2.740 11.480 3.000 ;
        RECT  10.470 2.230 10.730 3.000 ;
        RECT  9.510 2.740 10.470 3.000 ;
        RECT  9.250 2.280 9.510 3.000 ;
        RECT  7.375 2.740 9.250 3.000 ;
        RECT  7.215 2.245 7.375 3.000 ;
        RECT  2.810 2.740 7.215 3.000 ;
        RECT  2.550 2.570 2.810 3.000 ;
        RECT  0.690 2.740 2.550 3.000 ;
        RECT  0.690 1.810 0.930 1.970 ;
        RECT  0.530 1.810 0.690 3.000 ;
        RECT  0.000 2.740 0.530 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.695 1.190 10.970 1.450 ;
        RECT  10.485 0.615 10.695 1.890 ;
        RECT  10.155 0.615 10.485 0.895 ;
        RECT  10.105 1.730 10.485 1.890 ;
        RECT  10.045 1.345 10.305 1.550 ;
        RECT  9.845 1.730 10.105 2.305 ;
        RECT  8.850 1.380 10.045 1.550 ;
        RECT  9.035 1.730 9.845 1.890 ;
        RECT  8.690 0.665 8.850 2.175 ;
        RECT  7.715 2.400 8.815 2.560 ;
        RECT  8.475 0.665 8.690 0.890 ;
        RECT  8.355 1.915 8.690 2.175 ;
        RECT  8.055 0.685 8.115 1.555 ;
        RECT  7.955 0.685 8.055 2.145 ;
        RECT  7.895 1.330 7.955 2.145 ;
        RECT  6.895 1.330 7.895 1.555 ;
        RECT  7.555 1.735 7.715 2.560 ;
        RECT  6.555 1.735 7.555 1.895 ;
        RECT  6.215 2.075 7.035 2.235 ;
        RECT  6.735 1.295 6.895 1.555 ;
        RECT  6.395 0.650 6.555 1.895 ;
        RECT  5.120 0.650 6.395 0.810 ;
        RECT  6.055 0.990 6.215 2.235 ;
        RECT  5.805 1.995 6.055 2.235 ;
        RECT  5.645 1.995 5.805 2.560 ;
        RECT  5.460 1.040 5.695 1.200 ;
        RECT  3.390 2.400 5.645 2.560 ;
        RECT  5.300 1.040 5.460 2.220 ;
        RECT  3.730 2.060 5.300 2.220 ;
        RECT  4.960 0.650 5.120 1.880 ;
        RECT  4.925 0.650 4.960 0.810 ;
        RECT  4.515 1.720 4.960 1.880 ;
        RECT  4.345 0.880 4.605 1.140 ;
        RECT  4.085 0.880 4.345 1.040 ;
        RECT  3.925 0.705 4.085 1.040 ;
        RECT  3.635 0.880 3.925 1.040 ;
        RECT  3.570 2.015 3.730 2.220 ;
        RECT  3.635 1.675 3.700 1.835 ;
        RECT  3.475 0.880 3.635 1.835 ;
        RECT  2.385 2.015 3.570 2.175 ;
        RECT  3.440 1.675 3.475 1.835 ;
        RECT  3.130 2.355 3.390 2.560 ;
        RECT  2.725 0.610 2.955 0.870 ;
        RECT  2.565 0.325 2.725 0.870 ;
        RECT  1.235 0.325 2.565 0.485 ;
        RECT  2.380 2.015 2.385 2.380 ;
        RECT  2.220 0.665 2.380 2.380 ;
        RECT  1.855 0.665 2.220 0.825 ;
        RECT  1.575 2.220 2.220 2.380 ;
        RECT  1.880 1.035 2.040 2.035 ;
        RECT  1.465 1.035 1.880 1.195 ;
        RECT  1.305 0.925 1.465 1.195 ;
        RECT  0.815 0.925 1.305 1.085 ;
        RECT  0.975 0.325 1.235 0.585 ;
        RECT  0.555 0.785 0.815 1.085 ;
        RECT  0.285 0.925 0.555 1.085 ;
        RECT  0.285 2.200 0.335 2.460 ;
        RECT  0.125 0.925 0.285 2.460 ;
    END
END SDFFRQX1MTH

MACRO SDFFRQX2MTH
    CLASS CORE ;
    FOREIGN SDFFRQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.120 2.770 1.785 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.400 1.465 1.560 1.725 ;
        RECT  0.760 1.465 1.400 1.625 ;
        RECT  0.465 1.275 0.760 1.625 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 1.170 9.735 1.330 ;
        RECT  8.915 0.310 9.075 1.330 ;
        RECT  7.765 0.310 8.915 0.470 ;
        RECT  7.605 0.310 7.765 1.145 ;
        RECT  7.425 0.920 7.605 1.145 ;
        RECT  7.165 0.920 7.425 1.195 ;
        RECT  6.895 0.920 7.165 1.115 ;
        RECT  6.735 0.310 6.895 1.115 ;
        RECT  3.745 0.310 6.735 0.470 ;
        RECT  3.585 0.310 3.745 0.645 ;
        RECT  3.295 0.485 3.585 0.645 ;
        RECT  3.230 0.485 3.295 1.380 ;
        RECT  3.135 0.485 3.230 1.785 ;
        RECT  3.070 1.185 3.135 1.785 ;
        END
        AntennaGateArea 0.1664 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.170 0.375 11.380 2.410 ;
        RECT  11.095 0.375 11.170 0.975 ;
        RECT  11.095 1.810 11.170 2.410 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 2.150 1.220 2.545 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 1.330 4.450 1.540 ;
        RECT  3.830 1.220 3.990 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.815 -0.130 11.480 0.130 ;
        RECT  10.215 -0.130 10.815 0.335 ;
        RECT  9.965 -0.130 10.215 0.130 ;
        RECT  9.365 -0.130 9.965 0.355 ;
        RECT  7.425 -0.130 9.365 0.130 ;
        RECT  7.145 -0.130 7.425 0.740 ;
        RECT  3.405 -0.130 7.145 0.130 ;
        RECT  2.905 -0.130 3.405 0.300 ;
        RECT  0.725 -0.130 2.905 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.815 2.740 11.480 3.000 ;
        RECT  10.555 2.620 10.815 3.000 ;
        RECT  9.510 2.740 10.555 3.000 ;
        RECT  9.250 2.280 9.510 3.000 ;
        RECT  7.375 2.740 9.250 3.000 ;
        RECT  7.215 2.245 7.375 3.000 ;
        RECT  2.810 2.740 7.215 3.000 ;
        RECT  2.550 2.570 2.810 3.000 ;
        RECT  0.690 2.740 2.550 3.000 ;
        RECT  0.690 1.810 0.930 1.970 ;
        RECT  0.530 1.810 0.690 3.000 ;
        RECT  0.000 2.740 0.530 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.645 1.190 10.970 1.450 ;
        RECT  10.485 1.190 10.645 2.440 ;
        RECT  10.365 1.190 10.485 1.670 ;
        RECT  10.105 2.280 10.485 2.440 ;
        RECT  10.205 0.750 10.365 1.670 ;
        RECT  10.045 1.890 10.305 2.100 ;
        RECT  9.295 1.510 10.205 1.670 ;
        RECT  9.845 2.280 10.105 2.505 ;
        RECT  8.850 1.925 10.045 2.100 ;
        RECT  9.035 1.510 9.295 1.745 ;
        RECT  8.685 1.925 8.850 2.125 ;
        RECT  8.555 2.345 8.815 2.545 ;
        RECT  8.685 0.750 8.735 1.010 ;
        RECT  8.525 0.750 8.685 2.125 ;
        RECT  7.715 2.385 8.555 2.545 ;
        RECT  8.475 0.750 8.525 1.010 ;
        RECT  8.350 1.940 8.525 2.125 ;
        RECT  8.055 0.685 8.115 1.555 ;
        RECT  7.955 0.685 8.055 2.145 ;
        RECT  7.895 1.395 7.955 2.145 ;
        RECT  6.895 1.395 7.895 1.555 ;
        RECT  7.555 1.735 7.715 2.545 ;
        RECT  6.555 1.735 7.555 1.895 ;
        RECT  6.215 2.075 7.035 2.235 ;
        RECT  6.735 1.295 6.895 1.555 ;
        RECT  6.395 0.650 6.555 1.895 ;
        RECT  5.125 0.650 6.395 0.810 ;
        RECT  6.055 0.990 6.215 2.235 ;
        RECT  5.805 1.995 6.055 2.235 ;
        RECT  5.645 1.995 5.805 2.560 ;
        RECT  5.465 1.040 5.695 1.200 ;
        RECT  3.390 2.400 5.645 2.560 ;
        RECT  5.305 1.040 5.465 2.220 ;
        RECT  3.730 2.060 5.305 2.220 ;
        RECT  4.965 0.650 5.125 1.880 ;
        RECT  4.925 0.650 4.965 0.810 ;
        RECT  4.515 1.720 4.965 1.880 ;
        RECT  4.325 0.880 4.585 1.150 ;
        RECT  4.085 0.880 4.325 1.040 ;
        RECT  3.925 0.705 4.085 1.040 ;
        RECT  3.635 0.880 3.925 1.040 ;
        RECT  3.570 2.015 3.730 2.220 ;
        RECT  3.635 1.675 3.700 1.835 ;
        RECT  3.475 0.880 3.635 1.835 ;
        RECT  2.385 2.015 3.570 2.175 ;
        RECT  3.440 1.675 3.475 1.835 ;
        RECT  3.130 2.355 3.390 2.560 ;
        RECT  2.725 0.610 2.955 0.870 ;
        RECT  2.565 0.325 2.725 0.870 ;
        RECT  1.235 0.325 2.565 0.485 ;
        RECT  2.380 2.015 2.385 2.380 ;
        RECT  2.220 0.665 2.380 2.380 ;
        RECT  1.855 0.665 2.220 0.825 ;
        RECT  1.575 2.220 2.220 2.380 ;
        RECT  1.845 1.035 2.040 2.035 ;
        RECT  1.465 1.035 1.845 1.195 ;
        RECT  1.305 0.925 1.465 1.195 ;
        RECT  0.815 0.925 1.305 1.085 ;
        RECT  0.975 0.325 1.235 0.585 ;
        RECT  0.555 0.785 0.815 1.085 ;
        RECT  0.285 0.925 0.555 1.085 ;
        RECT  0.285 2.200 0.335 2.460 ;
        RECT  0.125 0.925 0.285 2.460 ;
    END
END SDFFRQX2MTH

MACRO SDFFRQX4MTH
    CLASS CORE ;
    FOREIGN SDFFRQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.120 2.770 1.785 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.400 1.465 1.560 1.725 ;
        RECT  0.760 1.465 1.400 1.625 ;
        RECT  0.465 1.275 0.760 1.625 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 1.170 9.735 1.330 ;
        RECT  8.915 0.310 9.075 1.330 ;
        RECT  7.765 0.310 8.915 0.470 ;
        RECT  7.605 0.310 7.765 1.145 ;
        RECT  7.165 0.920 7.605 1.145 ;
        RECT  6.895 0.920 7.165 1.115 ;
        RECT  6.735 0.310 6.895 1.115 ;
        RECT  3.745 0.310 6.735 0.470 ;
        RECT  3.585 0.310 3.745 0.645 ;
        RECT  3.295 0.485 3.585 0.645 ;
        RECT  3.230 0.485 3.295 1.380 ;
        RECT  3.135 0.485 3.230 1.785 ;
        RECT  3.070 1.185 3.135 1.785 ;
        END
        AntennaGateArea 0.2041 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.315 0.375 11.380 1.710 ;
        RECT  11.095 0.375 11.315 2.410 ;
        RECT  11.035 0.375 11.095 0.975 ;
        RECT  10.955 1.660 11.095 2.410 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 2.150 1.220 2.545 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  3.990 1.330 4.450 1.540 ;
        RECT  3.830 1.220 3.990 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.750 -0.130 11.890 0.130 ;
        RECT  10.490 -0.130 10.750 0.300 ;
        RECT  9.525 -0.130 10.490 0.130 ;
        RECT  9.265 -0.130 9.525 0.300 ;
        RECT  7.425 -0.130 9.265 0.130 ;
        RECT  7.145 -0.130 7.425 0.740 ;
        RECT  3.405 -0.130 7.145 0.130 ;
        RECT  2.905 -0.130 3.405 0.300 ;
        RECT  0.725 -0.130 2.905 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.755 2.740 11.890 3.000 ;
        RECT  11.495 1.890 11.755 3.000 ;
        RECT  10.675 2.740 11.495 3.000 ;
        RECT  10.415 2.620 10.675 3.000 ;
        RECT  9.510 2.740 10.415 3.000 ;
        RECT  9.250 2.280 9.510 3.000 ;
        RECT  7.375 2.740 9.250 3.000 ;
        RECT  7.215 2.245 7.375 3.000 ;
        RECT  2.810 2.740 7.215 3.000 ;
        RECT  2.550 2.570 2.810 3.000 ;
        RECT  0.690 2.740 2.550 3.000 ;
        RECT  0.690 1.810 0.930 1.970 ;
        RECT  0.530 1.810 0.690 3.000 ;
        RECT  0.000 2.740 0.530 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.645 1.220 10.915 1.480 ;
        RECT  10.485 1.220 10.645 2.440 ;
        RECT  10.385 1.220 10.485 1.670 ;
        RECT  10.105 2.280 10.485 2.440 ;
        RECT  10.120 0.750 10.385 1.670 ;
        RECT  10.045 1.890 10.305 2.100 ;
        RECT  9.295 1.510 10.120 1.670 ;
        RECT  9.845 2.280 10.105 2.515 ;
        RECT  8.850 1.925 10.045 2.100 ;
        RECT  9.035 1.510 9.295 1.745 ;
        RECT  8.685 1.925 8.850 2.125 ;
        RECT  7.715 2.385 8.815 2.545 ;
        RECT  8.685 0.750 8.735 1.010 ;
        RECT  8.525 0.750 8.685 2.125 ;
        RECT  8.475 0.750 8.525 1.010 ;
        RECT  8.350 1.940 8.525 2.125 ;
        RECT  8.055 0.685 8.115 1.555 ;
        RECT  7.955 0.685 8.055 2.145 ;
        RECT  7.895 1.395 7.955 2.145 ;
        RECT  6.895 1.395 7.895 1.555 ;
        RECT  7.555 1.735 7.715 2.545 ;
        RECT  6.555 1.735 7.555 1.895 ;
        RECT  6.215 2.075 7.035 2.235 ;
        RECT  6.735 1.295 6.895 1.555 ;
        RECT  6.395 0.650 6.555 1.895 ;
        RECT  5.120 0.650 6.395 0.810 ;
        RECT  6.055 0.990 6.215 2.235 ;
        RECT  5.805 1.995 6.055 2.235 ;
        RECT  5.645 1.995 5.805 2.560 ;
        RECT  5.460 1.040 5.695 1.200 ;
        RECT  3.390 2.400 5.645 2.560 ;
        RECT  5.300 1.040 5.460 2.220 ;
        RECT  3.730 2.060 5.300 2.220 ;
        RECT  4.960 0.650 5.120 1.880 ;
        RECT  4.925 0.650 4.960 0.810 ;
        RECT  4.515 1.720 4.960 1.880 ;
        RECT  4.345 0.880 4.605 1.150 ;
        RECT  4.085 0.880 4.345 1.040 ;
        RECT  3.925 0.705 4.085 1.040 ;
        RECT  3.635 0.880 3.925 1.040 ;
        RECT  3.570 2.015 3.730 2.220 ;
        RECT  3.635 1.675 3.700 1.835 ;
        RECT  3.475 0.880 3.635 1.835 ;
        RECT  2.385 2.015 3.570 2.175 ;
        RECT  3.440 1.675 3.475 1.835 ;
        RECT  3.130 2.355 3.390 2.560 ;
        RECT  2.720 0.610 2.955 0.870 ;
        RECT  2.560 0.325 2.720 0.870 ;
        RECT  1.235 0.325 2.560 0.485 ;
        RECT  2.380 2.015 2.385 2.380 ;
        RECT  2.220 0.665 2.380 2.380 ;
        RECT  1.855 0.665 2.220 0.825 ;
        RECT  1.575 2.220 2.220 2.380 ;
        RECT  1.845 1.035 2.040 2.035 ;
        RECT  1.465 1.035 1.845 1.195 ;
        RECT  1.305 0.925 1.465 1.195 ;
        RECT  0.815 0.925 1.305 1.085 ;
        RECT  0.975 0.325 1.235 0.585 ;
        RECT  0.555 0.795 0.815 1.085 ;
        RECT  0.285 0.925 0.555 1.085 ;
        RECT  0.285 2.200 0.335 2.460 ;
        RECT  0.125 0.925 0.285 2.460 ;
    END
END SDFFRQX4MTH

MACRO SDFFRX1MTH
    CLASS CORE ;
    FOREIGN SDFFRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.335 2.770 1.990 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 1.465 1.610 1.725 ;
        RECT  0.760 1.465 1.350 1.625 ;
        RECT  0.470 1.325 0.760 1.625 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.170 0.960 9.735 1.120 ;
        RECT  9.010 0.310 9.170 1.120 ;
        RECT  7.775 0.310 9.010 0.470 ;
        RECT  7.615 0.310 7.775 1.115 ;
        RECT  7.435 0.955 7.615 1.115 ;
        RECT  7.175 0.955 7.435 1.215 ;
        RECT  6.895 0.955 7.175 1.115 ;
        RECT  6.735 0.310 6.895 1.115 ;
        RECT  3.385 0.310 6.735 0.470 ;
        RECT  3.225 0.310 3.385 1.310 ;
        RECT  3.180 1.100 3.225 1.310 ;
        RECT  2.970 1.100 3.180 1.580 ;
        END
        AntennaGateArea 0.1586 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.765 1.290 10.970 1.580 ;
        RECT  10.735 1.290 10.765 1.995 ;
        RECT  10.575 0.815 10.735 1.995 ;
        END
        AntennaDiffArea 0.317 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.605 0.710 11.765 2.145 ;
        RECT  11.555 0.735 11.605 0.995 ;
        RECT  11.170 1.700 11.605 2.145 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 2.150 1.220 2.545 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 1.255 4.450 1.540 ;
        RECT  3.910 1.220 4.200 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.630 -0.130 11.890 0.130 ;
        RECT  10.690 -0.130 11.630 0.285 ;
        RECT  9.625 -0.130 10.690 0.130 ;
        RECT  9.365 -0.130 9.625 0.335 ;
        RECT  7.435 -0.130 9.365 0.130 ;
        RECT  7.275 -0.130 7.435 0.625 ;
        RECT  0.725 -0.130 7.275 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.530 2.740 11.890 3.000 ;
        RECT  10.270 2.545 10.530 3.000 ;
        RECT  9.365 2.740 10.270 3.000 ;
        RECT  9.105 2.360 9.365 3.000 ;
        RECT  7.375 2.740 9.105 3.000 ;
        RECT  7.215 2.245 7.375 3.000 ;
        RECT  2.880 2.740 7.215 3.000 ;
        RECT  2.620 2.560 2.880 3.000 ;
        RECT  0.690 2.740 2.620 3.000 ;
        RECT  0.690 1.810 0.930 1.970 ;
        RECT  0.515 1.810 0.690 3.000 ;
        RECT  0.000 2.740 0.515 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.360 1.240 11.415 1.500 ;
        RECT  11.200 0.470 11.360 1.500 ;
        RECT  10.415 0.470 11.200 0.630 ;
        RECT  10.395 0.355 10.415 0.630 ;
        RECT  10.235 0.355 10.395 2.005 ;
        RECT  10.155 0.355 10.235 0.515 ;
        RECT  9.950 1.845 10.235 2.005 ;
        RECT  9.895 1.300 10.055 1.650 ;
        RECT  9.690 1.845 9.950 2.535 ;
        RECT  8.635 1.300 9.895 1.460 ;
        RECT  9.295 1.845 9.690 2.005 ;
        RECT  9.035 1.640 9.295 2.005 ;
        RECT  7.715 2.385 8.815 2.545 ;
        RECT  8.635 0.705 8.735 0.865 ;
        RECT  8.475 0.705 8.635 2.185 ;
        RECT  8.355 1.925 8.475 2.185 ;
        RECT  7.955 0.655 8.115 2.145 ;
        RECT  7.895 1.395 7.955 2.145 ;
        RECT  6.905 1.395 7.895 1.555 ;
        RECT  7.555 1.735 7.715 2.545 ;
        RECT  6.555 1.735 7.555 1.895 ;
        RECT  6.215 2.075 7.035 2.235 ;
        RECT  6.745 1.295 6.905 1.555 ;
        RECT  6.395 0.650 6.555 1.895 ;
        RECT  5.120 0.650 6.395 0.810 ;
        RECT  6.055 0.990 6.215 2.235 ;
        RECT  5.810 1.995 6.055 2.235 ;
        RECT  5.650 1.995 5.810 2.560 ;
        RECT  5.470 1.040 5.695 1.200 ;
        RECT  3.550 2.400 5.650 2.560 ;
        RECT  5.310 1.040 5.470 2.220 ;
        RECT  4.185 2.060 5.310 2.220 ;
        RECT  4.960 0.650 5.120 1.880 ;
        RECT  4.860 0.650 4.960 0.825 ;
        RECT  4.520 1.720 4.960 1.880 ;
        RECT  4.425 0.880 4.685 1.075 ;
        RECT  4.005 0.880 4.425 1.040 ;
        RECT  4.025 2.015 4.185 2.220 ;
        RECT  3.110 2.015 4.025 2.175 ;
        RECT  3.745 0.650 4.005 1.040 ;
        RECT  3.725 1.675 3.790 1.835 ;
        RECT  3.725 0.880 3.745 1.040 ;
        RECT  3.565 0.880 3.725 1.835 ;
        RECT  3.530 1.675 3.565 1.835 ;
        RECT  3.290 2.355 3.550 2.560 ;
        RECT  2.950 2.015 3.110 2.380 ;
        RECT  2.885 0.325 3.045 0.920 ;
        RECT  2.380 2.220 2.950 2.380 ;
        RECT  1.325 0.325 2.885 0.485 ;
        RECT  2.220 0.665 2.380 2.380 ;
        RECT  1.945 0.665 2.220 0.825 ;
        RECT  1.575 2.220 2.220 2.380 ;
        RECT  1.880 1.035 2.040 2.035 ;
        RECT  1.465 1.035 1.880 1.195 ;
        RECT  1.305 0.985 1.465 1.195 ;
        RECT  1.165 0.325 1.325 0.805 ;
        RECT  0.815 0.985 1.305 1.145 ;
        RECT  1.065 0.645 1.165 0.805 ;
        RECT  0.555 0.765 0.815 1.145 ;
        RECT  0.285 0.985 0.555 1.145 ;
        RECT  0.285 2.165 0.335 2.425 ;
        RECT  0.125 0.985 0.285 2.425 ;
    END
END SDFFRX1MTH

MACRO SDFFRX2MTH
    CLASS CORE ;
    FOREIGN SDFFRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.300 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 0.880 2.770 1.710 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.350 1.465 1.610 1.725 ;
        RECT  0.760 1.465 1.350 1.625 ;
        RECT  0.465 1.325 0.760 1.625 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.210 1.040 9.890 1.200 ;
        RECT  9.050 0.325 9.210 1.200 ;
        RECT  7.845 0.325 9.050 0.485 ;
        RECT  7.685 0.325 7.845 1.115 ;
        RECT  6.895 0.955 7.685 1.115 ;
        RECT  6.735 0.310 6.895 1.115 ;
        RECT  3.385 0.310 6.735 0.470 ;
        RECT  3.225 0.310 3.385 1.535 ;
        RECT  3.180 1.050 3.225 1.535 ;
        RECT  2.970 1.050 3.180 1.580 ;
        END
        AntennaGateArea 0.169 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.180 1.290 11.380 1.580 ;
        RECT  11.030 0.815 11.180 2.285 ;
        RECT  11.020 0.765 11.030 2.285 ;
        RECT  10.870 0.765 11.020 1.025 ;
        RECT  10.840 1.685 11.020 2.285 ;
        END
        AntennaDiffArea 0.492 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.035 0.385 12.195 2.390 ;
        RECT  11.925 0.385 12.035 0.985 ;
        RECT  11.900 1.700 12.035 2.390 ;
        RECT  11.580 1.700 11.900 1.990 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 2.150 1.220 2.545 ;
        END
        AntennaGateArea 0.0715 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.200 1.330 4.450 1.540 ;
        RECT  3.970 1.220 4.200 1.540 ;
        RECT  3.905 1.220 3.970 1.505 ;
        END
        AntennaGateArea 0.0988 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.620 -0.130 12.300 0.130 ;
        RECT  11.360 -0.130 11.620 0.250 ;
        RECT  10.270 -0.130 11.360 0.130 ;
        RECT  10.010 -0.130 10.270 0.350 ;
        RECT  9.675 -0.130 10.010 0.130 ;
        RECT  9.415 -0.130 9.675 0.820 ;
        RECT  7.485 -0.130 9.415 0.130 ;
        RECT  7.225 -0.130 7.485 0.625 ;
        RECT  0.725 -0.130 7.225 0.130 ;
        RECT  0.125 -0.130 0.725 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.620 2.740 12.300 3.000 ;
        RECT  11.360 2.175 11.620 3.000 ;
        RECT  10.570 2.740 11.360 3.000 ;
        RECT  9.970 2.540 10.570 3.000 ;
        RECT  9.585 2.740 9.970 3.000 ;
        RECT  9.325 2.540 9.585 3.000 ;
        RECT  7.355 2.740 9.325 3.000 ;
        RECT  7.195 2.245 7.355 3.000 ;
        RECT  2.810 2.740 7.195 3.000 ;
        RECT  2.550 2.570 2.810 3.000 ;
        RECT  0.690 2.740 2.550 3.000 ;
        RECT  0.690 1.810 0.915 1.970 ;
        RECT  0.530 1.810 0.690 3.000 ;
        RECT  0.000 2.740 0.530 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.745 1.220 11.855 1.480 ;
        RECT  11.585 0.430 11.745 1.480 ;
        RECT  11.255 0.430 11.585 0.590 ;
        RECT  11.095 0.400 11.255 0.590 ;
        RECT  10.660 0.400 11.095 0.560 ;
        RECT  10.500 0.400 10.660 1.900 ;
        RECT  10.310 0.620 10.500 0.880 ;
        RECT  10.085 1.740 10.500 1.900 ;
        RECT  10.160 1.275 10.320 1.540 ;
        RECT  8.715 1.380 10.160 1.540 ;
        RECT  9.825 1.740 10.085 2.250 ;
        RECT  9.115 1.740 9.825 1.900 ;
        RECT  7.695 2.385 8.895 2.545 ;
        RECT  8.555 0.685 8.715 2.175 ;
        RECT  8.335 1.675 8.555 2.175 ;
        RECT  8.045 0.685 8.205 1.475 ;
        RECT  8.035 1.315 8.045 1.475 ;
        RECT  7.875 1.315 8.035 2.145 ;
        RECT  6.745 1.315 7.875 1.475 ;
        RECT  7.535 1.655 7.695 2.545 ;
        RECT  6.555 1.655 7.535 1.815 ;
        RECT  6.825 1.995 6.985 2.255 ;
        RECT  6.215 1.995 6.825 2.205 ;
        RECT  6.395 0.650 6.555 1.815 ;
        RECT  5.260 0.650 6.395 0.810 ;
        RECT  6.055 0.990 6.215 2.205 ;
        RECT  5.810 2.045 6.055 2.205 ;
        RECT  5.650 2.045 5.810 2.560 ;
        RECT  3.390 2.400 5.650 2.560 ;
        RECT  5.615 1.000 5.645 1.260 ;
        RECT  5.465 1.000 5.615 1.865 ;
        RECT  5.455 1.000 5.465 2.220 ;
        RECT  5.305 1.705 5.455 2.220 ;
        RECT  4.185 2.060 5.305 2.220 ;
        RECT  5.125 0.650 5.260 1.470 ;
        RECT  4.965 0.650 5.125 1.880 ;
        RECT  4.865 0.650 4.965 0.825 ;
        RECT  4.515 1.720 4.965 1.880 ;
        RECT  4.425 0.880 4.685 1.145 ;
        RECT  4.005 0.880 4.425 1.040 ;
        RECT  4.025 1.985 4.185 2.220 ;
        RECT  2.380 1.985 4.025 2.145 ;
        RECT  3.745 0.650 4.005 1.040 ;
        RECT  3.725 1.645 3.790 1.805 ;
        RECT  3.725 0.880 3.745 1.040 ;
        RECT  3.565 0.880 3.725 1.805 ;
        RECT  3.530 1.645 3.565 1.805 ;
        RECT  3.130 2.325 3.390 2.560 ;
        RECT  2.885 0.325 3.045 0.700 ;
        RECT  1.325 0.325 2.885 0.485 ;
        RECT  2.220 0.665 2.380 2.380 ;
        RECT  1.945 0.665 2.220 0.825 ;
        RECT  1.565 2.220 2.220 2.380 ;
        RECT  1.880 1.035 2.040 2.035 ;
        RECT  1.130 1.035 1.880 1.195 ;
        RECT  1.165 0.325 1.325 0.780 ;
        RECT  1.065 0.560 1.165 0.780 ;
        RECT  0.970 0.985 1.130 1.195 ;
        RECT  0.815 0.985 0.970 1.145 ;
        RECT  0.555 0.765 0.815 1.145 ;
        RECT  0.285 0.985 0.555 1.145 ;
        RECT  0.285 2.165 0.350 2.425 ;
        RECT  0.125 0.985 0.285 2.425 ;
    END
END SDFFRX2MTH

MACRO SDFFRX4MTH
    CLASS CORE ;
    FOREIGN SDFFRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.120 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.585 0.880 2.770 1.710 ;
        RECT  2.560 0.880 2.585 1.170 ;
        END
        AntennaGateArea 0.0689 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.540 1.465 1.630 1.715 ;
        RECT  1.330 1.110 1.540 1.715 ;
        RECT  0.625 1.110 1.330 1.270 ;
        RECT  0.465 0.985 0.625 1.270 ;
        END
        AntennaGateArea 0.1625 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.115 1.185 9.800 1.345 ;
        RECT  8.955 0.325 9.115 1.345 ;
        RECT  7.845 0.325 8.955 0.485 ;
        RECT  7.685 0.325 7.845 0.965 ;
        RECT  7.485 0.805 7.685 0.965 ;
        RECT  7.225 0.805 7.485 1.145 ;
        RECT  7.045 0.805 7.225 0.965 ;
        RECT  6.885 0.310 7.045 0.965 ;
        RECT  3.385 0.310 6.885 0.470 ;
        RECT  3.225 0.310 3.385 1.540 ;
        RECT  2.970 1.105 3.225 1.580 ;
        END
        AntennaGateArea 0.2301 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.200 0.815 11.460 2.285 ;
        RECT  11.145 0.815 11.200 0.975 ;
        RECT  11.170 1.290 11.200 1.580 ;
        END
        AntennaDiffArea 0.604 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.455 1.290 12.610 1.580 ;
        RECT  12.455 1.915 12.485 2.515 ;
        RECT  12.275 0.425 12.455 2.515 ;
        RECT  12.225 1.915 12.275 2.515 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.940 1.450 1.100 1.860 ;
        RECT  0.720 1.700 0.940 1.860 ;
        RECT  0.510 1.700 0.720 1.990 ;
        END
        AntennaGateArea 0.1417 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.255 4.450 1.540 ;
        RECT  3.905 1.255 4.160 1.515 ;
        END
        AntennaGateArea 0.1482 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.995 -0.130 13.120 0.130 ;
        RECT  12.735 -0.130 12.995 0.990 ;
        RECT  11.945 -0.130 12.735 0.130 ;
        RECT  11.685 -0.130 11.945 0.295 ;
        RECT  10.865 -0.130 11.685 0.130 ;
        RECT  10.605 -0.130 10.865 0.295 ;
        RECT  10.010 -0.130 10.605 0.130 ;
        RECT  9.410 -0.130 10.010 0.330 ;
        RECT  7.485 -0.130 9.410 0.130 ;
        RECT  7.225 -0.130 7.485 0.625 ;
        RECT  0.725 -0.130 7.225 0.130 ;
        RECT  0.125 -0.130 0.725 0.345 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.995 2.740 13.120 3.000 ;
        RECT  12.735 1.775 12.995 3.000 ;
        RECT  11.980 2.740 12.735 3.000 ;
        RECT  11.720 1.795 11.980 3.000 ;
        RECT  10.950 2.740 11.720 3.000 ;
        RECT  10.690 1.685 10.950 3.000 ;
        RECT  10.320 2.495 10.690 3.000 ;
        RECT  9.485 2.740 10.320 3.000 ;
        RECT  9.225 2.485 9.485 3.000 ;
        RECT  7.355 2.740 9.225 3.000 ;
        RECT  7.195 2.245 7.355 3.000 ;
        RECT  2.810 2.740 7.195 3.000 ;
        RECT  2.550 2.505 2.810 3.000 ;
        RECT  0.940 2.740 2.550 3.000 ;
        RECT  0.680 2.570 0.940 3.000 ;
        RECT  0.000 2.740 0.680 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.935 0.475 12.095 1.405 ;
        RECT  10.400 0.475 11.935 0.635 ;
        RECT  10.245 1.865 10.405 2.235 ;
        RECT  10.240 0.475 10.400 1.685 ;
        RECT  9.625 2.075 10.245 2.235 ;
        RECT  10.065 1.525 10.240 1.685 ;
        RECT  9.805 1.525 10.065 1.895 ;
        RECT  9.115 1.665 9.805 1.825 ;
        RECT  9.465 2.015 9.625 2.235 ;
        RECT  8.715 2.015 9.465 2.175 ;
        RECT  7.695 2.385 8.895 2.545 ;
        RECT  8.555 0.705 8.715 2.175 ;
        RECT  8.335 1.675 8.555 2.175 ;
        RECT  8.045 0.685 8.205 1.505 ;
        RECT  8.035 1.345 8.045 1.505 ;
        RECT  7.875 1.345 8.035 2.040 ;
        RECT  6.955 1.345 7.875 1.505 ;
        RECT  7.535 1.685 7.695 2.545 ;
        RECT  6.615 1.685 7.535 1.845 ;
        RECT  6.825 2.025 6.985 2.285 ;
        RECT  6.795 1.245 6.955 1.505 ;
        RECT  6.265 2.025 6.825 2.185 ;
        RECT  6.455 0.650 6.615 1.845 ;
        RECT  5.180 0.650 6.455 0.810 ;
        RECT  6.105 0.990 6.265 2.185 ;
        RECT  6.005 0.990 6.105 1.150 ;
        RECT  5.810 2.005 6.105 2.185 ;
        RECT  5.650 2.005 5.810 2.560 ;
        RECT  5.625 0.990 5.725 1.150 ;
        RECT  3.390 2.400 5.650 2.560 ;
        RECT  5.465 0.990 5.625 1.825 ;
        RECT  5.455 1.665 5.465 1.825 ;
        RECT  5.295 1.665 5.455 2.220 ;
        RECT  4.185 2.060 5.295 2.220 ;
        RECT  5.115 0.650 5.180 1.475 ;
        RECT  4.955 0.650 5.115 1.880 ;
        RECT  4.865 0.650 4.955 0.825 ;
        RECT  4.515 1.720 4.955 1.880 ;
        RECT  4.425 0.880 4.685 1.075 ;
        RECT  4.005 0.880 4.425 1.040 ;
        RECT  4.025 2.015 4.185 2.220 ;
        RECT  2.405 2.015 4.025 2.175 ;
        RECT  3.745 0.650 4.005 1.040 ;
        RECT  3.725 1.675 3.790 1.835 ;
        RECT  3.725 0.880 3.745 1.040 ;
        RECT  3.565 0.880 3.725 1.835 ;
        RECT  3.530 1.675 3.565 1.835 ;
        RECT  3.130 2.355 3.390 2.560 ;
        RECT  2.885 0.325 3.045 0.615 ;
        RECT  1.355 0.325 2.885 0.485 ;
        RECT  2.345 1.435 2.405 2.395 ;
        RECT  2.245 0.665 2.345 2.395 ;
        RECT  2.185 0.665 2.245 1.595 ;
        RECT  1.785 2.235 2.245 2.395 ;
        RECT  1.945 0.665 2.185 0.825 ;
        RECT  2.005 1.795 2.065 2.055 ;
        RECT  1.845 1.005 2.005 2.055 ;
        RECT  1.745 1.005 1.845 1.245 ;
        RECT  1.445 1.895 1.845 2.055 ;
        RECT  1.625 2.235 1.785 2.495 ;
        RECT  1.285 1.895 1.445 2.390 ;
        RECT  1.095 0.325 1.355 0.785 ;
        RECT  0.385 2.230 1.285 2.390 ;
        RECT  0.285 0.645 0.845 0.805 ;
        RECT  0.285 2.230 0.385 2.560 ;
        RECT  0.125 0.645 0.285 2.560 ;
    END
END SDFFRX4MTH

MACRO SDFFSHQX1MTH
    CLASS CORE ;
    FOREIGN SDFFSHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.585 1.100 6.950 1.705 ;
        END
        AntennaGateArea 0.1417 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.700 5.480 2.220 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.580 1.180 ;
        RECT  4.200 1.020 4.410 1.880 ;
        RECT  2.470 1.720 4.200 1.880 ;
        RECT  2.210 1.690 2.470 1.880 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.005 0.760 14.250 2.335 ;
        END
        AntennaDiffArea 0.34 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.845 3.680 1.170 ;
        RECT  3.380 0.845 3.540 1.520 ;
        END
        AntennaGateArea 0.0689 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.875 1.830 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.715 -0.130 14.350 0.130 ;
        RECT  13.505 -0.130 13.715 0.965 ;
        RECT  11.730 -0.130 13.505 0.130 ;
        RECT  11.470 -0.130 11.730 0.260 ;
        RECT  3.340 -0.130 11.470 0.130 ;
        RECT  3.180 -0.130 3.340 0.310 ;
        RECT  0.790 -0.130 3.180 0.130 ;
        RECT  0.290 -0.130 0.790 0.300 ;
        RECT  0.000 -0.130 0.290 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.745 2.740 14.350 3.000 ;
        RECT  13.505 1.735 13.745 3.000 ;
        RECT  12.915 2.570 13.505 3.000 ;
        RECT  10.170 2.740 12.915 3.000 ;
        RECT  9.910 2.620 10.170 3.000 ;
        RECT  9.000 2.740 9.910 3.000 ;
        RECT  8.740 2.620 9.000 3.000 ;
        RECT  6.600 2.740 8.740 3.000 ;
        RECT  6.000 2.620 6.600 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.325 1.220 13.695 1.480 ;
        RECT  13.165 0.370 13.325 2.335 ;
        RECT  12.595 0.370 13.165 0.530 ;
        RECT  12.490 2.175 13.165 2.335 ;
        RECT  12.825 0.765 12.985 1.995 ;
        RECT  12.775 1.205 12.825 1.995 ;
        RECT  12.495 1.205 12.775 1.470 ;
        RECT  12.335 0.310 12.595 0.530 ;
        RECT  12.330 2.175 12.490 2.455 ;
        RECT  12.315 0.775 12.475 0.935 ;
        RECT  12.035 0.370 12.335 0.530 ;
        RECT  11.270 2.295 12.330 2.455 ;
        RECT  12.155 0.775 12.315 1.775 ;
        RECT  12.070 1.515 12.155 1.775 ;
        RECT  11.910 1.515 12.070 2.115 ;
        RECT  11.875 0.370 12.035 0.635 ;
        RECT  11.390 1.955 11.910 2.115 ;
        RECT  11.170 0.475 11.875 0.635 ;
        RECT  11.570 0.815 11.730 1.775 ;
        RECT  10.830 0.815 11.570 0.975 ;
        RECT  11.230 1.155 11.390 2.115 ;
        RECT  10.490 1.155 11.230 1.315 ;
        RECT  11.010 0.375 11.170 0.635 ;
        RECT  10.890 1.495 11.050 2.440 ;
        RECT  9.550 2.270 10.890 2.440 ;
        RECT  10.670 0.310 10.830 0.975 ;
        RECT  10.610 1.920 10.710 2.080 ;
        RECT  3.680 0.310 10.670 0.470 ;
        RECT  10.450 1.575 10.610 2.080 ;
        RECT  10.330 0.650 10.490 1.315 ;
        RECT  10.150 1.575 10.450 1.735 ;
        RECT  6.360 0.650 10.330 0.810 ;
        RECT  9.990 0.990 10.150 1.735 ;
        RECT  9.890 0.990 9.990 1.150 ;
        RECT  9.230 1.575 9.990 1.735 ;
        RECT  8.420 1.915 9.750 2.075 ;
        RECT  9.450 0.990 9.710 1.395 ;
        RECT  9.290 2.270 9.550 2.500 ;
        RECT  8.420 0.990 9.450 1.150 ;
        RECT  8.440 2.270 9.290 2.440 ;
        RECT  8.970 1.330 9.230 1.735 ;
        RECT  8.280 2.270 8.440 2.470 ;
        RECT  8.260 0.990 8.420 2.075 ;
        RECT  7.760 2.300 8.280 2.470 ;
        RECT  8.100 1.840 8.260 2.075 ;
        RECT  7.940 1.840 8.100 2.120 ;
        RECT  7.760 1.005 7.840 1.325 ;
        RECT  7.600 1.005 7.760 2.470 ;
        RECT  5.820 2.280 7.600 2.440 ;
        RECT  7.260 1.485 7.420 2.100 ;
        RECT  5.920 1.940 7.260 2.100 ;
        RECT  6.200 0.650 6.360 1.760 ;
        RECT  6.100 1.600 6.200 1.760 ;
        RECT  5.760 0.650 5.920 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.210 0.650 5.760 0.810 ;
        RECT  4.750 1.360 5.760 1.520 ;
        RECT  1.665 2.400 5.660 2.560 ;
        RECT  4.020 0.650 4.900 0.810 ;
        RECT  2.005 2.060 4.840 2.220 ;
        RECT  4.590 1.360 4.750 1.870 ;
        RECT  3.860 0.650 4.020 1.540 ;
        RECT  3.720 1.380 3.860 1.540 ;
        RECT  3.520 0.310 3.680 0.665 ;
        RECT  2.955 0.505 3.520 0.665 ;
        RECT  2.795 0.505 2.955 1.540 ;
        RECT  2.750 0.505 2.795 0.665 ;
        RECT  2.695 1.260 2.795 1.540 ;
        RECT  2.590 0.365 2.750 0.665 ;
        RECT  2.110 1.260 2.695 1.420 ;
        RECT  1.130 0.310 2.410 0.470 ;
        RECT  1.950 1.160 2.110 1.420 ;
        RECT  1.845 1.860 2.005 2.220 ;
        RECT  1.770 1.860 1.845 2.020 ;
        RECT  1.610 0.650 1.770 2.020 ;
        RECT  1.505 2.200 1.665 2.560 ;
        RECT  1.310 0.650 1.610 0.810 ;
        RECT  1.430 2.200 1.505 2.360 ;
        RECT  1.270 1.110 1.430 2.360 ;
        RECT  0.970 0.310 1.130 0.930 ;
        RECT  0.385 0.770 0.970 0.930 ;
        RECT  0.285 0.770 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.770 0.285 2.290 ;
    END
END SDFFSHQX1MTH

MACRO SDFFSHQX2MTH
    CLASS CORE ;
    FOREIGN SDFFSHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.760 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.585 1.100 6.950 1.710 ;
        END
        AntennaGateArea 0.1677 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.700 5.480 2.220 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.580 1.180 ;
        RECT  4.200 1.020 4.410 1.880 ;
        RECT  2.470 1.720 4.200 1.880 ;
        RECT  2.210 1.690 2.470 1.880 ;
        END
        AntennaGateArea 0.1313 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.375 0.400 14.660 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.845 3.680 1.170 ;
        RECT  3.380 0.845 3.540 1.520 ;
        END
        AntennaGateArea 0.0988 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.760 1.830 ;
        END
        AntennaGateArea 0.1508 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.125 -0.130 14.760 0.130 ;
        RECT  13.915 -0.130 14.125 0.955 ;
        RECT  12.140 -0.130 13.915 0.130 ;
        RECT  11.880 -0.130 12.140 0.260 ;
        RECT  3.340 -0.130 11.880 0.130 ;
        RECT  3.180 -0.130 3.340 0.310 ;
        RECT  0.790 -0.130 3.180 0.130 ;
        RECT  0.290 -0.130 0.790 0.300 ;
        RECT  0.000 -0.130 0.290 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.945 2.740 14.760 3.000 ;
        RECT  13.305 2.570 13.945 3.000 ;
        RECT  9.930 2.740 13.305 3.000 ;
        RECT  9.670 2.620 9.930 3.000 ;
        RECT  9.010 2.740 9.670 3.000 ;
        RECT  8.750 2.620 9.010 3.000 ;
        RECT  6.600 2.740 8.750 3.000 ;
        RECT  6.000 2.620 6.600 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.915 1.185 14.100 1.445 ;
        RECT  13.755 1.185 13.915 2.335 ;
        RECT  13.735 1.185 13.755 1.445 ;
        RECT  13.035 2.175 13.755 2.335 ;
        RECT  13.575 0.370 13.735 1.445 ;
        RECT  13.180 0.370 13.575 0.530 ;
        RECT  13.390 1.735 13.490 1.995 ;
        RECT  13.230 0.815 13.390 1.995 ;
        RECT  13.115 1.205 13.230 1.470 ;
        RECT  12.865 0.310 13.180 0.530 ;
        RECT  12.875 2.175 13.035 2.455 ;
        RECT  12.800 0.775 12.915 0.935 ;
        RECT  11.910 2.295 12.875 2.455 ;
        RECT  12.445 0.370 12.865 0.530 ;
        RECT  12.660 0.775 12.800 1.775 ;
        RECT  12.610 0.775 12.660 2.115 ;
        RECT  12.500 1.515 12.610 2.115 ;
        RECT  11.980 1.955 12.500 2.115 ;
        RECT  12.285 0.370 12.445 0.600 ;
        RECT  12.160 0.780 12.320 1.775 ;
        RECT  11.310 0.440 12.285 0.600 ;
        RECT  11.130 0.780 12.160 0.940 ;
        RECT  11.820 1.120 11.980 2.115 ;
        RECT  10.790 1.120 11.820 1.280 ;
        RECT  11.465 1.460 11.625 2.430 ;
        RECT  11.080 1.460 11.465 1.620 ;
        RECT  9.500 2.270 11.465 2.430 ;
        RECT  10.310 1.910 11.285 2.070 ;
        RECT  10.970 0.310 11.130 0.940 ;
        RECT  3.680 0.310 10.970 0.470 ;
        RECT  10.630 0.650 10.790 1.280 ;
        RECT  6.360 0.650 10.630 0.810 ;
        RECT  10.310 0.990 10.430 1.150 ;
        RECT  10.150 0.990 10.310 2.070 ;
        RECT  10.000 1.585 10.150 2.070 ;
        RECT  9.230 1.585 10.000 1.745 ;
        RECT  9.660 0.990 9.920 1.405 ;
        RECT  8.260 1.925 9.750 2.085 ;
        RECT  8.260 0.990 9.660 1.150 ;
        RECT  9.340 2.270 9.500 2.550 ;
        RECT  8.440 2.270 9.340 2.430 ;
        RECT  8.970 1.330 9.230 1.745 ;
        RECT  8.280 2.270 8.440 2.470 ;
        RECT  7.760 2.300 8.280 2.470 ;
        RECT  8.100 0.990 8.260 2.085 ;
        RECT  7.940 1.840 8.100 2.120 ;
        RECT  7.760 1.065 7.840 1.335 ;
        RECT  7.600 1.065 7.760 2.470 ;
        RECT  5.820 2.280 7.600 2.440 ;
        RECT  7.260 1.485 7.420 2.100 ;
        RECT  5.920 1.940 7.260 2.100 ;
        RECT  6.200 0.650 6.360 1.760 ;
        RECT  6.100 1.600 6.200 1.760 ;
        RECT  5.760 0.650 5.920 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.210 0.650 5.760 0.810 ;
        RECT  4.750 1.360 5.760 1.520 ;
        RECT  1.665 2.400 5.660 2.560 ;
        RECT  4.020 0.650 4.900 0.810 ;
        RECT  2.005 2.060 4.840 2.220 ;
        RECT  4.590 1.360 4.750 1.870 ;
        RECT  3.860 0.650 4.020 1.540 ;
        RECT  3.750 1.380 3.860 1.540 ;
        RECT  3.520 0.310 3.680 0.665 ;
        RECT  2.785 0.505 3.520 0.665 ;
        RECT  2.770 1.260 2.955 1.540 ;
        RECT  2.770 0.385 2.785 0.665 ;
        RECT  2.695 0.385 2.770 1.540 ;
        RECT  2.610 0.385 2.695 1.420 ;
        RECT  2.110 1.260 2.610 1.420 ;
        RECT  1.130 0.310 2.430 0.470 ;
        RECT  1.950 1.160 2.110 1.420 ;
        RECT  1.845 1.860 2.005 2.220 ;
        RECT  1.770 1.860 1.845 2.020 ;
        RECT  1.610 0.650 1.770 2.020 ;
        RECT  1.505 2.200 1.665 2.560 ;
        RECT  1.310 0.650 1.610 0.810 ;
        RECT  1.430 2.200 1.505 2.360 ;
        RECT  1.270 1.110 1.430 2.360 ;
        RECT  0.970 0.310 1.130 0.930 ;
        RECT  0.385 0.770 0.970 0.930 ;
        RECT  0.285 0.770 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.770 0.285 2.290 ;
    END
END SDFFSHQX2MTH

MACRO SDFFSHQX4MTH
    CLASS CORE ;
    FOREIGN SDFFSHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.170 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.640 1.100 6.950 1.705 ;
        END
        AntennaGateArea 0.1989 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.270 2.060 5.480 2.220 ;
        RECT  5.020 1.700 5.270 2.220 ;
        END
        AntennaGateArea 0.0611 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.550 1.180 ;
        RECT  4.200 1.020 4.410 1.880 ;
        RECT  2.405 1.720 4.200 1.880 ;
        RECT  2.145 1.690 2.405 1.880 ;
        END
        AntennaGateArea 0.1781 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.575 1.285 14.660 1.595 ;
        RECT  14.320 0.400 14.575 2.370 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.880 3.680 1.170 ;
        RECT  3.380 0.880 3.540 1.520 ;
        END
        AntennaGateArea 0.1417 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.760 1.830 ;
        END
        AntennaGateArea 0.1833 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.995 -0.130 15.170 0.130 ;
        RECT  14.835 -0.130 14.995 1.000 ;
        RECT  13.995 -0.130 14.835 0.130 ;
        RECT  13.395 -0.130 13.995 0.250 ;
        RECT  12.140 -0.130 13.395 0.130 ;
        RECT  11.880 -0.130 12.140 0.260 ;
        RECT  3.120 -0.130 11.880 0.130 ;
        RECT  2.860 -0.130 3.120 0.250 ;
        RECT  0.700 -0.130 2.860 0.130 ;
        RECT  0.200 -0.130 0.700 0.365 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.995 2.740 15.170 3.000 ;
        RECT  14.835 1.810 14.995 3.000 ;
        RECT  13.945 2.740 14.835 3.000 ;
        RECT  13.305 2.570 13.945 3.000 ;
        RECT  8.980 2.740 13.305 3.000 ;
        RECT  8.720 2.620 8.980 3.000 ;
        RECT  6.600 2.740 8.720 3.000 ;
        RECT  6.000 2.620 6.600 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.915 1.215 14.115 1.475 ;
        RECT  13.755 0.465 13.915 2.335 ;
        RECT  13.155 0.465 13.755 0.625 ;
        RECT  13.615 1.215 13.755 1.475 ;
        RECT  13.115 2.175 13.755 2.335 ;
        RECT  13.405 1.735 13.505 1.995 ;
        RECT  13.245 0.815 13.405 1.995 ;
        RECT  13.135 1.215 13.245 1.475 ;
        RECT  12.995 0.370 13.155 0.625 ;
        RECT  12.955 2.175 13.115 2.465 ;
        RECT  12.445 0.370 12.995 0.565 ;
        RECT  11.910 2.305 12.955 2.465 ;
        RECT  12.770 1.525 12.865 1.785 ;
        RECT  12.770 0.785 12.825 0.945 ;
        RECT  12.605 0.785 12.770 2.125 ;
        RECT  12.565 0.785 12.605 0.945 ;
        RECT  11.995 1.965 12.605 2.125 ;
        RECT  12.285 0.370 12.445 0.635 ;
        RECT  12.175 0.815 12.335 1.785 ;
        RECT  11.520 0.475 12.285 0.635 ;
        RECT  10.830 0.815 12.175 0.975 ;
        RECT  11.835 1.155 11.995 2.125 ;
        RECT  10.490 1.155 11.835 1.315 ;
        RECT  11.465 1.495 11.625 2.435 ;
        RECT  11.020 0.375 11.520 0.635 ;
        RECT  11.040 1.495 11.465 1.655 ;
        RECT  9.550 2.275 11.465 2.435 ;
        RECT  10.150 1.930 11.285 2.090 ;
        RECT  10.670 0.310 10.830 0.975 ;
        RECT  3.645 0.310 10.670 0.470 ;
        RECT  10.330 0.650 10.490 1.315 ;
        RECT  6.440 0.650 10.330 0.810 ;
        RECT  9.990 0.990 10.150 2.090 ;
        RECT  9.890 0.990 9.990 1.150 ;
        RECT  9.230 1.595 9.990 1.755 ;
        RECT  8.260 1.935 9.750 2.095 ;
        RECT  9.450 0.990 9.710 1.415 ;
        RECT  9.290 2.275 9.550 2.500 ;
        RECT  8.260 0.990 9.450 1.150 ;
        RECT  8.440 2.275 9.290 2.435 ;
        RECT  8.970 1.330 9.230 1.755 ;
        RECT  8.280 2.275 8.440 2.475 ;
        RECT  7.740 2.305 8.280 2.475 ;
        RECT  8.100 0.990 8.260 2.095 ;
        RECT  8.080 1.840 8.100 2.095 ;
        RECT  7.920 1.840 8.080 2.120 ;
        RECT  7.740 1.180 7.840 1.440 ;
        RECT  7.580 1.180 7.740 2.475 ;
        RECT  5.820 2.280 7.580 2.440 ;
        RECT  7.240 1.660 7.400 2.100 ;
        RECT  5.890 1.940 7.240 2.100 ;
        RECT  6.280 0.650 6.440 1.760 ;
        RECT  6.070 1.600 6.280 1.760 ;
        RECT  5.730 0.650 5.890 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.150 0.650 5.730 0.810 ;
        RECT  4.750 1.360 5.730 1.520 ;
        RECT  1.615 2.400 5.660 2.560 ;
        RECT  4.020 0.650 4.900 0.810 ;
        RECT  1.955 2.060 4.840 2.220 ;
        RECT  4.590 1.360 4.750 1.870 ;
        RECT  3.860 0.650 4.020 1.540 ;
        RECT  3.720 1.380 3.860 1.540 ;
        RECT  3.485 0.310 3.645 0.665 ;
        RECT  2.905 0.505 3.485 0.665 ;
        RECT  2.905 1.260 2.955 1.540 ;
        RECT  2.745 0.505 2.905 1.540 ;
        RECT  2.530 0.505 2.745 0.665 ;
        RECT  2.695 1.260 2.745 1.540 ;
        RECT  2.080 1.260 2.695 1.420 ;
        RECT  2.370 0.385 2.530 0.665 ;
        RECT  1.040 0.310 2.160 0.470 ;
        RECT  1.920 1.160 2.080 1.420 ;
        RECT  1.795 1.675 1.955 2.220 ;
        RECT  1.740 1.675 1.795 1.835 ;
        RECT  1.580 0.650 1.740 1.835 ;
        RECT  1.455 2.200 1.615 2.560 ;
        RECT  1.220 0.650 1.580 0.810 ;
        RECT  1.400 2.200 1.455 2.360 ;
        RECT  1.240 1.110 1.400 2.360 ;
        RECT  0.880 0.310 1.040 0.930 ;
        RECT  0.385 0.770 0.880 0.930 ;
        RECT  0.285 0.770 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.770 0.285 2.290 ;
    END
END SDFFSHQX4MTH

MACRO SDFFSHQX8MTH
    CLASS CORE ;
    FOREIGN SDFFSHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.640 1.100 6.950 1.705 ;
        END
        AntennaGateArea 0.2002 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.270 2.060 5.480 2.220 ;
        RECT  5.020 1.700 5.270 2.220 ;
        END
        AntennaGateArea 0.0611 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.550 1.180 ;
        RECT  4.200 1.020 4.410 1.880 ;
        RECT  2.405 1.720 4.200 1.880 ;
        RECT  2.145 1.690 2.405 1.880 ;
        END
        AntennaGateArea 0.1781 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.505 0.400 15.765 2.370 ;
        RECT  14.760 1.285 15.505 1.595 ;
        RECT  14.465 0.400 14.760 2.410 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 0.880 3.680 1.170 ;
        RECT  3.380 0.880 3.540 1.520 ;
        END
        AntennaGateArea 0.1417 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.760 1.830 ;
        END
        AntennaGateArea 0.1833 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.275 -0.130 16.400 0.130 ;
        RECT  16.015 -0.130 16.275 1.000 ;
        RECT  15.255 -0.130 16.015 0.130 ;
        RECT  14.995 -0.130 15.255 1.000 ;
        RECT  14.285 -0.130 14.995 0.130 ;
        RECT  14.025 -0.130 14.285 1.000 ;
        RECT  13.605 -0.130 14.025 0.250 ;
        RECT  12.140 -0.130 13.605 0.130 ;
        RECT  11.880 -0.130 12.140 0.260 ;
        RECT  3.120 -0.130 11.880 0.130 ;
        RECT  2.860 -0.130 3.120 0.250 ;
        RECT  0.700 -0.130 2.860 0.130 ;
        RECT  0.200 -0.130 0.700 0.375 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.275 2.740 16.400 3.000 ;
        RECT  16.015 1.805 16.275 3.000 ;
        RECT  15.255 2.740 16.015 3.000 ;
        RECT  14.995 1.805 15.255 3.000 ;
        RECT  14.285 2.740 14.995 3.000 ;
        RECT  14.025 1.805 14.285 3.000 ;
        RECT  13.300 2.570 14.025 3.000 ;
        RECT  9.010 2.740 13.300 3.000 ;
        RECT  8.750 2.620 9.010 3.000 ;
        RECT  6.600 2.740 8.750 3.000 ;
        RECT  6.000 2.620 6.600 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.845 1.215 14.215 1.475 ;
        RECT  13.685 0.465 13.845 2.335 ;
        RECT  13.225 0.465 13.685 0.625 ;
        RECT  13.115 2.175 13.685 2.335 ;
        RECT  13.405 0.815 13.505 0.975 ;
        RECT  13.405 1.685 13.505 1.945 ;
        RECT  13.245 0.815 13.405 1.945 ;
        RECT  13.135 1.215 13.245 1.475 ;
        RECT  13.065 0.370 13.225 0.625 ;
        RECT  12.955 2.175 13.115 2.465 ;
        RECT  12.445 0.370 13.065 0.565 ;
        RECT  11.910 2.305 12.955 2.465 ;
        RECT  12.770 1.525 12.865 1.785 ;
        RECT  12.770 0.785 12.825 0.945 ;
        RECT  12.605 0.785 12.770 2.125 ;
        RECT  12.565 0.785 12.605 0.945 ;
        RECT  11.995 1.965 12.605 2.125 ;
        RECT  12.285 0.370 12.445 0.635 ;
        RECT  12.175 0.815 12.335 1.785 ;
        RECT  11.520 0.475 12.285 0.635 ;
        RECT  10.830 0.815 12.175 0.975 ;
        RECT  11.835 1.155 11.995 2.125 ;
        RECT  10.490 1.155 11.835 1.315 ;
        RECT  11.465 1.495 11.625 2.435 ;
        RECT  11.020 0.375 11.520 0.635 ;
        RECT  11.040 1.495 11.465 1.655 ;
        RECT  9.550 2.275 11.465 2.435 ;
        RECT  10.150 1.930 11.285 2.090 ;
        RECT  10.670 0.310 10.830 0.975 ;
        RECT  3.645 0.310 10.670 0.470 ;
        RECT  10.330 0.650 10.490 1.315 ;
        RECT  6.440 0.650 10.330 0.810 ;
        RECT  9.990 0.990 10.150 2.090 ;
        RECT  9.890 0.990 9.990 1.150 ;
        RECT  9.230 1.595 9.990 1.755 ;
        RECT  8.260 1.935 9.750 2.095 ;
        RECT  9.450 0.990 9.710 1.415 ;
        RECT  9.290 2.275 9.550 2.500 ;
        RECT  8.260 0.990 9.450 1.150 ;
        RECT  8.440 2.275 9.290 2.435 ;
        RECT  8.970 1.330 9.230 1.755 ;
        RECT  8.280 2.275 8.440 2.470 ;
        RECT  7.740 2.305 8.280 2.470 ;
        RECT  8.100 0.990 8.260 2.095 ;
        RECT  8.080 1.840 8.100 2.095 ;
        RECT  7.920 1.840 8.080 2.120 ;
        RECT  7.740 1.180 7.840 1.440 ;
        RECT  7.580 1.180 7.740 2.470 ;
        RECT  5.820 2.280 7.580 2.440 ;
        RECT  7.240 1.660 7.400 2.100 ;
        RECT  5.890 1.940 7.240 2.100 ;
        RECT  6.280 0.650 6.440 1.760 ;
        RECT  6.070 1.600 6.280 1.760 ;
        RECT  5.730 0.650 5.890 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.150 0.650 5.730 0.810 ;
        RECT  4.750 1.360 5.730 1.520 ;
        RECT  1.615 2.400 5.660 2.560 ;
        RECT  4.020 0.650 4.900 0.810 ;
        RECT  1.955 2.060 4.840 2.220 ;
        RECT  4.590 1.360 4.750 1.870 ;
        RECT  3.860 0.650 4.020 1.540 ;
        RECT  3.720 1.380 3.860 1.540 ;
        RECT  3.485 0.310 3.645 0.665 ;
        RECT  2.905 0.505 3.485 0.665 ;
        RECT  2.905 1.260 2.955 1.540 ;
        RECT  2.745 0.505 2.905 1.540 ;
        RECT  2.530 0.505 2.745 0.665 ;
        RECT  2.695 1.260 2.745 1.540 ;
        RECT  2.080 1.260 2.695 1.420 ;
        RECT  2.370 0.385 2.530 0.665 ;
        RECT  1.040 0.310 2.160 0.470 ;
        RECT  1.920 1.160 2.080 1.420 ;
        RECT  1.795 1.675 1.955 2.220 ;
        RECT  1.740 1.675 1.795 1.835 ;
        RECT  1.580 0.650 1.740 1.835 ;
        RECT  1.455 2.200 1.615 2.560 ;
        RECT  1.220 0.650 1.580 0.810 ;
        RECT  1.400 2.200 1.455 2.360 ;
        RECT  1.240 1.110 1.400 2.360 ;
        RECT  0.880 0.310 1.040 0.930 ;
        RECT  0.385 0.770 0.880 0.930 ;
        RECT  0.285 0.770 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.770 0.285 2.290 ;
    END
END SDFFSHQX8MTH

MACRO SDFFSQX1MTH
    CLASS CORE ;
    FOREIGN SDFFSQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.370 1.330 9.470 1.490 ;
        RECT  9.080 1.330 9.370 1.540 ;
        RECT  8.765 1.380 9.080 1.540 ;
        RECT  8.605 1.380 8.765 2.560 ;
        RECT  8.205 2.400 8.605 2.560 ;
        END
        AntennaGateArea 0.1079 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.260 1.650 1.520 ;
        RECT  0.920 1.260 1.560 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.035 0.360 1.755 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 1.700 10.970 2.055 ;
        RECT  10.785 0.760 10.945 2.055 ;
        RECT  10.735 0.760 10.785 1.020 ;
        RECT  10.685 1.700 10.785 2.055 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 1.045 2.265 1.305 ;
        RECT  1.990 1.145 2.105 1.305 ;
        RECT  1.830 1.145 1.990 2.055 ;
        RECT  1.740 1.700 1.830 2.055 ;
        RECT  1.315 1.895 1.740 2.055 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.320 4.815 1.480 ;
        RECT  4.025 1.320 4.450 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 -0.130 11.070 0.130 ;
        RECT  10.145 -0.130 10.405 0.250 ;
        RECT  9.815 -0.130 10.145 0.130 ;
        RECT  9.215 -0.130 9.815 0.250 ;
        RECT  4.445 -0.130 9.215 0.130 ;
        RECT  4.185 -0.130 4.445 0.250 ;
        RECT  0.675 -0.130 4.185 0.130 ;
        RECT  0.175 -0.130 0.675 0.300 ;
        RECT  0.000 -0.130 0.175 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 2.740 11.070 3.000 ;
        RECT  9.805 2.570 10.405 3.000 ;
        RECT  9.525 2.740 9.805 3.000 ;
        RECT  9.265 2.570 9.525 3.000 ;
        RECT  8.025 2.740 9.265 3.000 ;
        RECT  7.425 2.620 8.025 3.000 ;
        RECT  7.235 2.740 7.425 3.000 ;
        RECT  6.635 2.620 7.235 3.000 ;
        RECT  5.790 2.740 6.635 3.000 ;
        RECT  5.630 2.570 5.790 3.000 ;
        RECT  0.385 2.740 5.630 3.000 ;
        RECT  0.125 2.230 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.370 1.190 10.605 1.450 ;
        RECT  10.210 0.605 10.370 2.180 ;
        RECT  9.720 0.605 10.210 0.765 ;
        RECT  9.160 2.020 10.210 2.180 ;
        RECT  9.930 1.265 10.030 1.525 ;
        RECT  9.770 0.990 9.930 1.525 ;
        RECT  7.995 0.990 9.770 1.150 ;
        RECT  8.945 2.020 9.160 2.320 ;
        RECT  8.835 0.605 8.935 0.765 ;
        RECT  8.675 0.310 8.835 0.765 ;
        RECT  5.525 0.310 8.675 0.470 ;
        RECT  7.995 1.880 8.420 2.145 ;
        RECT  7.835 0.765 7.995 2.440 ;
        RECT  6.840 2.280 7.835 2.440 ;
        RECT  7.425 0.650 7.475 0.975 ;
        RECT  7.335 1.910 7.460 2.070 ;
        RECT  7.335 0.650 7.425 1.025 ;
        RECT  7.175 0.650 7.335 2.070 ;
        RECT  6.315 0.650 7.175 0.810 ;
        RECT  6.785 0.990 6.945 1.570 ;
        RECT  6.680 1.990 6.840 2.440 ;
        RECT  6.625 0.990 6.785 1.520 ;
        RECT  6.380 1.360 6.625 1.520 ;
        RECT  6.285 1.360 6.380 2.250 ;
        RECT  6.265 0.650 6.315 0.965 ;
        RECT  6.220 1.360 6.285 2.390 ;
        RECT  6.105 0.650 6.265 1.015 ;
        RECT  6.120 1.990 6.220 2.390 ;
        RECT  5.450 2.230 6.120 2.390 ;
        RECT  5.425 0.800 6.105 0.965 ;
        RECT  5.865 1.190 6.025 1.450 ;
        RECT  5.770 1.290 5.865 1.450 ;
        RECT  5.610 1.290 5.770 1.880 ;
        RECT  4.885 1.720 5.610 1.880 ;
        RECT  5.265 0.310 5.525 0.620 ;
        RECT  5.290 2.230 5.450 2.560 ;
        RECT  5.265 0.800 5.425 1.540 ;
        RECT  2.710 2.400 5.290 2.560 ;
        RECT  4.335 0.800 5.265 0.965 ;
        RECT  5.135 1.380 5.265 1.540 ;
        RECT  3.290 2.060 5.110 2.220 ;
        RECT  3.840 0.430 5.020 0.590 ;
        RECT  4.625 1.690 4.885 1.880 ;
        RECT  3.825 1.720 4.625 1.880 ;
        RECT  4.175 0.800 4.335 1.140 ;
        RECT  4.075 0.980 4.175 1.140 ;
        RECT  3.825 0.310 3.840 0.590 ;
        RECT  3.665 0.310 3.825 1.880 ;
        RECT  3.575 0.310 3.665 0.590 ;
        RECT  3.470 1.520 3.665 1.780 ;
        RECT  3.325 0.770 3.485 1.030 ;
        RECT  3.290 0.870 3.325 1.030 ;
        RECT  3.130 0.870 3.290 2.220 ;
        RECT  2.785 0.365 2.945 2.220 ;
        RECT  1.275 0.365 2.785 0.525 ;
        RECT  2.525 2.060 2.785 2.220 ;
        RECT  2.445 0.705 2.605 1.645 ;
        RECT  2.365 2.060 2.525 2.475 ;
        RECT  1.650 0.705 2.445 0.865 ;
        RECT  2.330 1.485 2.445 1.645 ;
        RECT  0.925 2.315 2.365 2.475 ;
        RECT  2.170 1.485 2.330 1.785 ;
        RECT  1.490 0.705 1.650 0.985 ;
        RECT  0.815 0.825 1.490 0.985 ;
        RECT  1.115 0.335 1.275 0.595 ;
        RECT  0.665 2.215 0.925 2.475 ;
        RECT  0.700 0.765 0.815 1.025 ;
        RECT  0.700 1.755 0.815 1.915 ;
        RECT  0.540 0.765 0.700 1.915 ;
    END
END SDFFSQX1MTH

MACRO SDFFSQX2MTH
    CLASS CORE ;
    FOREIGN SDFFSQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.370 1.330 9.470 1.490 ;
        RECT  9.080 1.330 9.370 1.540 ;
        RECT  8.765 1.380 9.080 1.540 ;
        RECT  8.605 1.380 8.765 2.560 ;
        RECT  8.205 2.400 8.605 2.560 ;
        END
        AntennaGateArea 0.1092 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.260 1.650 1.520 ;
        RECT  0.920 1.260 1.560 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.035 0.360 1.755 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 1.700 10.970 1.990 ;
        RECT  10.785 0.400 10.945 2.390 ;
        RECT  10.685 0.400 10.785 1.000 ;
        RECT  10.760 1.700 10.785 2.390 ;
        RECT  10.685 1.790 10.760 2.390 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 1.045 2.265 1.305 ;
        RECT  1.990 1.145 2.105 1.305 ;
        RECT  1.830 1.145 1.990 2.055 ;
        RECT  1.740 1.700 1.830 2.055 ;
        RECT  1.315 1.895 1.740 2.055 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.320 4.815 1.480 ;
        RECT  4.025 1.320 4.450 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 -0.130 11.070 0.130 ;
        RECT  10.145 -0.130 10.405 0.250 ;
        RECT  9.815 -0.130 10.145 0.130 ;
        RECT  9.215 -0.130 9.815 0.250 ;
        RECT  4.445 -0.130 9.215 0.130 ;
        RECT  4.185 -0.130 4.445 0.250 ;
        RECT  0.675 -0.130 4.185 0.130 ;
        RECT  0.175 -0.130 0.675 0.300 ;
        RECT  0.000 -0.130 0.175 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.405 2.740 11.070 3.000 ;
        RECT  9.805 2.570 10.405 3.000 ;
        RECT  9.525 2.740 9.805 3.000 ;
        RECT  9.265 2.570 9.525 3.000 ;
        RECT  8.025 2.740 9.265 3.000 ;
        RECT  7.425 2.620 8.025 3.000 ;
        RECT  7.235 2.740 7.425 3.000 ;
        RECT  6.635 2.620 7.235 3.000 ;
        RECT  5.790 2.740 6.635 3.000 ;
        RECT  5.630 2.570 5.790 3.000 ;
        RECT  0.385 2.740 5.630 3.000 ;
        RECT  0.125 2.230 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.370 1.190 10.605 1.450 ;
        RECT  10.210 0.605 10.370 2.180 ;
        RECT  9.720 0.605 10.210 0.765 ;
        RECT  9.105 2.020 10.210 2.180 ;
        RECT  9.930 1.265 10.030 1.525 ;
        RECT  9.770 0.990 9.930 1.525 ;
        RECT  7.995 0.990 9.770 1.150 ;
        RECT  8.945 2.020 9.105 2.355 ;
        RECT  8.835 0.605 8.935 0.765 ;
        RECT  8.675 0.310 8.835 0.765 ;
        RECT  5.525 0.310 8.675 0.470 ;
        RECT  7.995 1.880 8.420 2.145 ;
        RECT  7.835 0.765 7.995 2.440 ;
        RECT  6.840 2.280 7.835 2.440 ;
        RECT  7.425 0.650 7.475 0.975 ;
        RECT  7.335 1.910 7.460 2.070 ;
        RECT  7.335 0.650 7.425 1.025 ;
        RECT  7.175 0.650 7.335 2.070 ;
        RECT  6.265 0.650 7.175 0.810 ;
        RECT  6.945 1.360 6.995 1.520 ;
        RECT  6.885 1.310 6.945 1.570 ;
        RECT  6.785 0.990 6.885 1.570 ;
        RECT  6.680 1.990 6.840 2.440 ;
        RECT  6.625 0.990 6.785 1.520 ;
        RECT  6.380 1.360 6.625 1.520 ;
        RECT  6.285 1.360 6.380 2.250 ;
        RECT  6.220 1.360 6.285 2.390 ;
        RECT  6.105 0.650 6.265 1.015 ;
        RECT  6.120 1.990 6.220 2.390 ;
        RECT  5.450 2.230 6.120 2.390 ;
        RECT  5.425 0.800 6.105 0.965 ;
        RECT  5.865 1.190 6.025 1.450 ;
        RECT  5.770 1.290 5.865 1.450 ;
        RECT  5.610 1.290 5.770 1.880 ;
        RECT  4.885 1.720 5.610 1.880 ;
        RECT  5.265 0.310 5.525 0.620 ;
        RECT  5.290 2.230 5.450 2.560 ;
        RECT  5.265 0.800 5.425 1.540 ;
        RECT  2.710 2.400 5.290 2.560 ;
        RECT  4.335 0.800 5.265 0.965 ;
        RECT  5.135 1.380 5.265 1.540 ;
        RECT  3.290 2.060 5.110 2.220 ;
        RECT  3.840 0.430 5.020 0.590 ;
        RECT  4.625 1.690 4.885 1.880 ;
        RECT  3.825 1.720 4.625 1.880 ;
        RECT  4.175 0.800 4.335 1.140 ;
        RECT  4.075 0.980 4.175 1.140 ;
        RECT  3.825 0.310 3.840 0.590 ;
        RECT  3.665 0.310 3.825 1.880 ;
        RECT  3.575 0.310 3.665 0.590 ;
        RECT  3.470 1.520 3.665 1.780 ;
        RECT  3.325 0.770 3.485 1.030 ;
        RECT  3.290 0.870 3.325 1.030 ;
        RECT  3.130 0.870 3.290 2.220 ;
        RECT  2.785 0.365 2.945 2.220 ;
        RECT  1.275 0.365 2.785 0.525 ;
        RECT  2.525 2.060 2.785 2.220 ;
        RECT  2.445 0.705 2.605 1.645 ;
        RECT  2.365 2.060 2.525 2.475 ;
        RECT  1.650 0.705 2.445 0.865 ;
        RECT  2.330 1.485 2.445 1.645 ;
        RECT  0.925 2.315 2.365 2.475 ;
        RECT  2.170 1.485 2.330 1.785 ;
        RECT  1.490 0.705 1.650 0.985 ;
        RECT  0.815 0.825 1.490 0.985 ;
        RECT  1.115 0.335 1.275 0.595 ;
        RECT  0.665 2.215 0.925 2.475 ;
        RECT  0.700 0.765 0.815 1.025 ;
        RECT  0.700 1.755 0.815 1.915 ;
        RECT  0.540 0.765 0.700 1.915 ;
    END
END SDFFSQX2MTH

MACRO SDFFSQX4MTH
    CLASS CORE ;
    FOREIGN SDFFSQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.370 1.330 9.470 1.490 ;
        RECT  9.080 1.330 9.370 1.540 ;
        RECT  8.765 1.380 9.080 1.540 ;
        RECT  8.605 1.380 8.765 2.560 ;
        RECT  8.205 2.400 8.605 2.560 ;
        END
        AntennaGateArea 0.1092 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.560 1.260 1.650 1.520 ;
        RECT  0.920 1.260 1.560 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.035 0.360 1.755 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 1.700 10.970 1.990 ;
        RECT  10.890 1.700 10.945 2.390 ;
        RECT  10.680 0.400 10.890 2.390 ;
        RECT  10.650 1.790 10.680 2.390 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.105 1.045 2.265 1.305 ;
        RECT  1.990 1.145 2.105 1.305 ;
        RECT  1.830 1.145 1.990 2.055 ;
        RECT  1.740 1.700 1.830 2.055 ;
        RECT  1.315 1.895 1.740 2.055 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.320 4.815 1.480 ;
        RECT  4.025 1.320 4.450 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.350 -0.130 11.480 0.130 ;
        RECT  10.090 -0.130 10.350 0.295 ;
        RECT  9.815 -0.130 10.090 0.130 ;
        RECT  9.215 -0.130 9.815 0.250 ;
        RECT  4.445 -0.130 9.215 0.130 ;
        RECT  4.185 -0.130 4.445 0.250 ;
        RECT  0.675 -0.130 4.185 0.130 ;
        RECT  0.175 -0.130 0.675 0.300 ;
        RECT  0.000 -0.130 0.175 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.270 2.740 11.480 3.000 ;
        RECT  9.770 2.570 10.270 3.000 ;
        RECT  9.525 2.740 9.770 3.000 ;
        RECT  9.265 2.570 9.525 3.000 ;
        RECT  8.025 2.740 9.265 3.000 ;
        RECT  7.425 2.620 8.025 3.000 ;
        RECT  7.235 2.740 7.425 3.000 ;
        RECT  6.635 2.620 7.235 3.000 ;
        RECT  5.790 2.740 6.635 3.000 ;
        RECT  5.630 2.570 5.790 3.000 ;
        RECT  0.385 2.740 5.630 3.000 ;
        RECT  0.125 2.230 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.370 1.190 10.500 1.450 ;
        RECT  10.210 0.615 10.370 2.180 ;
        RECT  9.720 0.615 10.210 0.775 ;
        RECT  9.105 2.020 10.210 2.180 ;
        RECT  9.930 1.265 10.030 1.525 ;
        RECT  9.770 0.990 9.930 1.525 ;
        RECT  7.995 0.990 9.770 1.150 ;
        RECT  8.945 2.020 9.105 2.355 ;
        RECT  8.835 0.605 8.935 0.765 ;
        RECT  8.675 0.310 8.835 0.765 ;
        RECT  5.525 0.310 8.675 0.470 ;
        RECT  7.995 1.880 8.420 2.145 ;
        RECT  7.835 0.765 7.995 2.440 ;
        RECT  6.840 2.280 7.835 2.440 ;
        RECT  7.335 1.910 7.460 2.070 ;
        RECT  7.335 0.650 7.425 1.025 ;
        RECT  7.175 0.650 7.335 2.070 ;
        RECT  6.265 0.650 7.175 0.810 ;
        RECT  6.625 0.990 6.945 1.570 ;
        RECT  6.680 1.990 6.840 2.440 ;
        RECT  6.380 1.375 6.625 1.570 ;
        RECT  6.285 1.375 6.380 2.250 ;
        RECT  6.220 1.375 6.285 2.390 ;
        RECT  6.105 0.650 6.265 1.015 ;
        RECT  6.120 1.990 6.220 2.390 ;
        RECT  5.450 2.230 6.120 2.390 ;
        RECT  5.425 0.810 6.105 0.975 ;
        RECT  5.865 1.190 6.025 1.450 ;
        RECT  5.770 1.290 5.865 1.450 ;
        RECT  5.610 1.290 5.770 1.880 ;
        RECT  4.885 1.720 5.610 1.880 ;
        RECT  5.265 0.310 5.525 0.620 ;
        RECT  5.290 2.230 5.450 2.560 ;
        RECT  5.265 0.810 5.425 1.540 ;
        RECT  2.710 2.400 5.290 2.560 ;
        RECT  4.335 0.810 5.265 0.975 ;
        RECT  5.135 1.380 5.265 1.540 ;
        RECT  3.290 2.060 5.110 2.220 ;
        RECT  4.755 0.360 5.020 0.590 ;
        RECT  4.625 1.690 4.885 1.880 ;
        RECT  3.840 0.430 4.755 0.590 ;
        RECT  3.825 1.720 4.625 1.880 ;
        RECT  4.175 0.810 4.335 1.140 ;
        RECT  4.075 0.980 4.175 1.140 ;
        RECT  3.825 0.310 3.840 0.590 ;
        RECT  3.665 0.310 3.825 1.880 ;
        RECT  3.575 0.310 3.665 0.590 ;
        RECT  3.470 1.520 3.665 1.780 ;
        RECT  3.325 0.770 3.485 1.030 ;
        RECT  3.290 0.870 3.325 1.030 ;
        RECT  3.130 0.870 3.290 2.220 ;
        RECT  2.785 0.365 2.945 2.220 ;
        RECT  1.275 0.365 2.785 0.525 ;
        RECT  2.525 2.060 2.785 2.220 ;
        RECT  2.445 0.705 2.605 1.645 ;
        RECT  2.365 2.060 2.525 2.475 ;
        RECT  1.650 0.705 2.445 0.865 ;
        RECT  2.330 1.485 2.445 1.645 ;
        RECT  0.925 2.315 2.365 2.475 ;
        RECT  2.170 1.485 2.330 1.785 ;
        RECT  1.490 0.705 1.650 0.985 ;
        RECT  0.815 0.825 1.490 0.985 ;
        RECT  1.115 0.335 1.275 0.595 ;
        RECT  0.665 2.215 0.925 2.475 ;
        RECT  0.700 0.765 0.815 1.025 ;
        RECT  0.700 1.755 0.815 1.915 ;
        RECT  0.540 0.765 0.700 1.915 ;
    END
END SDFFSQX4MTH

MACRO SDFFSRHQX1MTH
    CLASS CORE ;
    FOREIGN SDFFSRHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.540 1.045 6.870 1.660 ;
        END
        AntennaGateArea 0.1365 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.700 5.480 2.220 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.540 1.180 ;
        RECT  4.250 1.020 4.410 1.880 ;
        RECT  4.160 1.290 4.250 1.880 ;
        RECT  2.420 1.720 4.160 1.880 ;
        RECT  2.255 1.620 2.420 1.880 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.640 1.385 12.900 1.590 ;
        RECT  10.600 1.430 12.640 1.590 ;
        RECT  10.310 1.330 10.600 1.590 ;
        END
        AntennaGateArea 0.1391 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.090 0.765 16.300 2.115 ;
        RECT  16.015 0.765 16.090 1.025 ;
        RECT  16.015 1.850 16.090 2.115 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.065 0.845 3.640 1.170 ;
        END
        AntennaGateArea 0.0598 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.760 1.830 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.175 -0.130 16.400 0.130 ;
        RECT  15.575 -0.130 16.175 0.255 ;
        RECT  15.355 -0.130 15.575 0.130 ;
        RECT  14.415 -0.130 15.355 0.255 ;
        RECT  3.385 -0.130 14.415 0.130 ;
        RECT  3.125 -0.130 3.385 0.310 ;
        RECT  0.830 -0.130 3.125 0.130 ;
        RECT  0.330 -0.130 0.830 0.300 ;
        RECT  0.000 -0.130 0.330 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.680 2.740 16.400 3.000 ;
        RECT  15.080 2.570 15.680 3.000 ;
        RECT  10.860 2.740 15.080 3.000 ;
        RECT  10.600 2.620 10.860 3.000 ;
        RECT  9.920 2.740 10.600 3.000 ;
        RECT  9.660 2.620 9.920 3.000 ;
        RECT  8.800 2.740 9.660 3.000 ;
        RECT  8.540 2.620 8.800 3.000 ;
        RECT  6.930 2.740 8.540 3.000 ;
        RECT  5.990 2.620 6.930 3.000 ;
        RECT  0.815 2.740 5.990 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.580 1.205 15.910 1.465 ;
        RECT  15.420 0.435 15.580 2.285 ;
        RECT  14.020 0.435 15.420 0.595 ;
        RECT  15.310 1.205 15.420 1.465 ;
        RECT  14.825 2.125 15.420 2.285 ;
        RECT  15.100 1.685 15.240 1.945 ;
        RECT  15.100 0.815 15.195 0.975 ;
        RECT  14.935 0.815 15.100 1.945 ;
        RECT  14.870 1.255 14.935 1.515 ;
        RECT  14.665 2.125 14.825 2.515 ;
        RECT  12.790 2.355 14.665 2.515 ;
        RECT  14.405 1.625 14.550 1.885 ;
        RECT  14.405 0.885 14.455 1.045 ;
        RECT  14.245 0.885 14.405 2.175 ;
        RECT  14.195 0.885 14.245 1.045 ;
        RECT  13.240 2.015 14.245 2.175 ;
        RECT  13.680 1.675 14.050 1.835 ;
        RECT  13.860 0.355 14.020 0.725 ;
        RECT  12.100 0.355 13.860 0.515 ;
        RECT  13.520 0.695 13.680 1.835 ;
        RECT  11.920 0.695 13.520 0.855 ;
        RECT  13.080 1.035 13.240 2.175 ;
        RECT  11.580 1.035 13.080 1.195 ;
        RECT  12.760 1.865 13.080 2.025 ;
        RECT  12.530 2.295 12.790 2.515 ;
        RECT  11.470 1.815 12.250 1.975 ;
        RECT  11.730 2.185 11.990 2.440 ;
        RECT  11.760 0.310 11.920 0.855 ;
        RECT  3.730 0.310 11.760 0.470 ;
        RECT  9.360 2.270 11.730 2.440 ;
        RECT  11.420 0.650 11.580 1.195 ;
        RECT  11.310 1.815 11.470 2.090 ;
        RECT  6.320 0.650 11.420 0.810 ;
        RECT  9.850 1.930 11.310 2.090 ;
        RECT  11.080 0.990 11.240 1.250 ;
        RECT  9.850 0.990 11.080 1.150 ;
        RECT  9.690 0.990 9.850 2.090 ;
        RECT  9.600 1.470 9.690 1.730 ;
        RECT  9.240 0.990 9.460 1.250 ;
        RECT  9.100 2.270 9.360 2.560 ;
        RECT  9.080 0.990 9.240 2.090 ;
        RECT  8.230 2.270 9.100 2.440 ;
        RECT  8.900 1.840 9.080 2.090 ;
        RECT  8.260 1.840 8.900 2.000 ;
        RECT  8.260 0.990 8.480 1.150 ;
        RECT  8.100 0.990 8.260 2.000 ;
        RECT  8.070 2.270 8.230 2.500 ;
        RECT  7.890 1.840 8.100 2.000 ;
        RECT  7.550 2.300 8.070 2.500 ;
        RECT  7.730 1.840 7.890 2.120 ;
        RECT  7.550 1.005 7.800 1.265 ;
        RECT  7.390 1.005 7.550 2.500 ;
        RECT  5.820 2.280 7.390 2.440 ;
        RECT  7.050 1.325 7.210 2.100 ;
        RECT  5.880 1.940 7.050 2.100 ;
        RECT  6.160 0.650 6.320 1.760 ;
        RECT  6.060 1.600 6.160 1.760 ;
        RECT  5.720 0.650 5.880 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.170 0.650 5.720 0.810 ;
        RECT  4.750 1.360 5.720 1.520 ;
        RECT  1.665 2.400 5.660 2.560 ;
        RECT  4.070 0.650 4.860 0.810 ;
        RECT  2.005 2.060 4.820 2.220 ;
        RECT  4.590 1.360 4.750 1.870 ;
        RECT  3.980 0.650 4.070 1.110 ;
        RECT  3.910 0.650 3.980 1.540 ;
        RECT  3.820 0.950 3.910 1.540 ;
        RECT  3.720 1.380 3.820 1.540 ;
        RECT  3.570 0.310 3.730 0.665 ;
        RECT  2.855 0.505 3.570 0.665 ;
        RECT  2.855 1.380 2.955 1.540 ;
        RECT  2.725 0.505 2.855 1.540 ;
        RECT  2.695 0.365 2.725 1.540 ;
        RECT  2.565 0.365 2.695 1.295 ;
        RECT  2.110 1.135 2.565 1.295 ;
        RECT  1.170 0.310 2.385 0.470 ;
        RECT  1.950 1.135 2.110 1.400 ;
        RECT  1.845 1.860 2.005 2.220 ;
        RECT  1.770 1.860 1.845 2.020 ;
        RECT  1.610 0.650 1.770 2.020 ;
        RECT  1.505 2.200 1.665 2.560 ;
        RECT  1.350 0.650 1.610 0.810 ;
        RECT  1.100 2.200 1.505 2.360 ;
        RECT  1.270 1.110 1.430 1.370 ;
        RECT  1.100 1.210 1.270 1.370 ;
        RECT  1.010 0.310 1.170 0.925 ;
        RECT  0.940 1.210 1.100 2.360 ;
        RECT  0.385 0.765 1.010 0.925 ;
        RECT  0.285 0.765 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.765 0.285 2.290 ;
    END
END SDFFSRHQX1MTH

MACRO SDFFSRHQX2MTH
    CLASS CORE ;
    FOREIGN SDFFSRHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.810 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 1.020 6.990 1.660 ;
        END
        AntennaGateArea 0.1599 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.020 1.700 5.480 2.220 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.580 1.180 ;
        RECT  4.250 1.020 4.410 1.880 ;
        RECT  4.140 1.265 4.250 1.880 ;
        RECT  2.565 1.720 4.140 1.880 ;
        RECT  2.305 1.665 2.565 1.880 ;
        END
        AntennaGateArea 0.1066 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.055 1.385 13.315 1.635 ;
        RECT  11.790 1.475 13.055 1.635 ;
        RECT  11.530 1.440 11.790 1.635 ;
        RECT  11.010 1.475 11.530 1.635 ;
        RECT  10.720 1.330 11.010 1.635 ;
        RECT  10.580 1.440 10.720 1.635 ;
        END
        AntennaGateArea 0.1677 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.500 0.400 16.710 2.405 ;
        RECT  16.425 0.400 16.500 1.000 ;
        RECT  16.425 1.685 16.500 2.405 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.590 0.845 3.620 1.105 ;
        RECT  3.380 0.845 3.590 1.520 ;
        END
        AntennaGateArea 0.0858 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.760 1.830 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.200 -0.130 16.810 0.130 ;
        RECT  15.940 -0.130 16.200 0.955 ;
        RECT  15.385 -0.130 15.940 0.130 ;
        RECT  14.785 -0.130 15.385 0.260 ;
        RECT  3.390 -0.130 14.785 0.130 ;
        RECT  3.230 -0.130 3.390 0.310 ;
        RECT  0.795 -0.130 3.230 0.130 ;
        RECT  0.295 -0.130 0.795 0.300 ;
        RECT  0.000 -0.130 0.295 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.030 2.740 16.810 3.000 ;
        RECT  15.430 2.570 16.030 3.000 ;
        RECT  11.100 2.740 15.430 3.000 ;
        RECT  10.840 2.620 11.100 3.000 ;
        RECT  10.160 2.740 10.840 3.000 ;
        RECT  9.900 2.620 10.160 3.000 ;
        RECT  9.010 2.740 9.900 3.000 ;
        RECT  8.750 2.620 9.010 3.000 ;
        RECT  7.420 2.740 8.750 3.000 ;
        RECT  6.820 2.620 7.420 3.000 ;
        RECT  6.600 2.740 6.820 3.000 ;
        RECT  6.000 2.620 6.600 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.920 1.205 16.100 1.465 ;
        RECT  15.760 1.205 15.920 2.235 ;
        RECT  15.600 0.475 15.760 1.465 ;
        RECT  15.110 2.075 15.760 2.235 ;
        RECT  14.445 0.475 15.600 0.635 ;
        RECT  15.270 1.735 15.580 1.895 ;
        RECT  15.270 0.815 15.420 0.975 ;
        RECT  15.110 0.815 15.270 1.895 ;
        RECT  15.000 1.140 15.110 1.400 ;
        RECT  14.950 2.075 15.110 2.455 ;
        RECT  14.375 2.295 14.950 2.455 ;
        RECT  14.750 1.625 14.840 1.885 ;
        RECT  14.590 0.825 14.750 2.115 ;
        RECT  14.395 0.825 14.590 0.985 ;
        RECT  13.655 1.955 14.590 2.115 ;
        RECT  14.185 0.355 14.445 0.635 ;
        RECT  13.995 1.615 14.410 1.775 ;
        RECT  14.110 2.295 14.375 2.515 ;
        RECT  12.430 0.355 14.185 0.515 ;
        RECT  12.820 2.295 14.110 2.455 ;
        RECT  13.835 0.695 13.995 1.775 ;
        RECT  12.250 0.695 13.835 0.855 ;
        RECT  13.495 1.035 13.655 2.115 ;
        RECT  11.910 1.035 13.495 1.195 ;
        RECT  13.050 1.865 13.495 2.115 ;
        RECT  12.280 1.815 12.540 2.005 ;
        RECT  11.780 1.845 12.280 2.005 ;
        RECT  12.020 2.185 12.280 2.440 ;
        RECT  12.090 0.310 12.250 0.855 ;
        RECT  3.730 0.310 12.090 0.470 ;
        RECT  9.570 2.270 12.020 2.440 ;
        RECT  11.750 0.650 11.910 1.195 ;
        RECT  11.620 1.845 11.780 2.090 ;
        RECT  6.360 0.650 11.750 0.810 ;
        RECT  10.290 1.930 11.620 2.090 ;
        RECT  11.410 0.990 11.570 1.250 ;
        RECT  10.290 0.990 11.410 1.150 ;
        RECT  10.130 0.990 10.290 2.090 ;
        RECT  9.900 0.990 10.130 1.150 ;
        RECT  9.840 1.455 10.130 1.715 ;
        RECT  9.310 2.270 9.570 2.560 ;
        RECT  9.380 1.015 9.550 1.340 ;
        RECT  9.220 1.015 9.380 2.090 ;
        RECT  8.440 2.270 9.310 2.440 ;
        RECT  9.110 1.840 9.220 2.090 ;
        RECT  8.260 1.840 9.110 2.000 ;
        RECT  8.260 0.990 8.520 1.150 ;
        RECT  8.280 2.270 8.440 2.480 ;
        RECT  7.760 2.300 8.280 2.480 ;
        RECT  8.100 0.990 8.260 2.000 ;
        RECT  7.940 1.840 8.100 2.120 ;
        RECT  7.760 1.005 7.840 1.275 ;
        RECT  7.600 1.005 7.760 2.480 ;
        RECT  5.820 2.280 7.600 2.440 ;
        RECT  7.260 1.485 7.420 2.100 ;
        RECT  5.920 1.940 7.260 2.100 ;
        RECT  6.200 0.650 6.360 1.760 ;
        RECT  6.100 1.600 6.200 1.760 ;
        RECT  5.760 0.650 5.920 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.210 0.650 5.760 0.810 ;
        RECT  4.750 1.360 5.760 1.520 ;
        RECT  1.665 2.400 5.660 2.560 ;
        RECT  4.070 0.650 4.900 0.810 ;
        RECT  2.005 2.060 4.840 2.220 ;
        RECT  4.590 1.360 4.750 1.870 ;
        RECT  3.960 0.650 4.070 1.055 ;
        RECT  3.910 0.650 3.960 1.540 ;
        RECT  3.800 0.845 3.910 1.540 ;
        RECT  3.770 1.280 3.800 1.540 ;
        RECT  3.570 0.310 3.730 0.665 ;
        RECT  2.855 0.505 3.570 0.665 ;
        RECT  2.855 1.380 2.955 1.540 ;
        RECT  2.695 0.395 2.855 1.540 ;
        RECT  2.615 0.395 2.695 1.300 ;
        RECT  2.205 1.140 2.615 1.300 ;
        RECT  1.135 0.310 2.435 0.470 ;
        RECT  2.045 1.085 2.205 1.345 ;
        RECT  1.865 1.860 2.005 2.220 ;
        RECT  1.845 0.650 1.865 2.220 ;
        RECT  1.705 0.650 1.845 2.020 ;
        RECT  1.315 0.650 1.705 0.810 ;
        RECT  1.505 2.200 1.665 2.560 ;
        RECT  1.365 1.110 1.525 1.370 ;
        RECT  1.100 2.200 1.505 2.360 ;
        RECT  1.100 1.210 1.365 1.370 ;
        RECT  0.975 0.310 1.135 0.790 ;
        RECT  0.940 1.210 1.100 2.360 ;
        RECT  0.385 0.630 0.975 0.790 ;
        RECT  0.285 0.630 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.630 0.285 2.290 ;
    END
END SDFFSRHQX2MTH

MACRO SDFFSRHQX4MTH
    CLASS CORE ;
    FOREIGN SDFFSRHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.220 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.655 1.150 6.990 1.750 ;
        END
        AntennaGateArea 0.1807 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.270 2.060 5.480 2.220 ;
        RECT  5.020 1.700 5.270 2.220 ;
        END
        AntennaGateArea 0.0715 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.580 1.180 ;
        RECT  4.360 1.020 4.410 1.580 ;
        RECT  4.250 1.020 4.360 1.880 ;
        RECT  4.200 1.250 4.250 1.880 ;
        RECT  2.420 1.720 4.200 1.880 ;
        RECT  2.260 1.620 2.420 1.880 ;
        END
        AntennaGateArea 0.1287 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.910 1.385 13.315 1.545 ;
        RECT  11.750 1.385 11.910 1.635 ;
        RECT  11.010 1.475 11.750 1.635 ;
        RECT  10.720 1.330 11.010 1.635 ;
        RECT  10.540 1.440 10.720 1.635 ;
        END
        AntennaGateArea 0.2041 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.585 1.290 16.715 1.580 ;
        RECT  16.325 0.400 16.585 2.400 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 0.875 3.640 1.200 ;
        END
        AntennaGateArea 0.13 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.510 1.235 0.800 1.830 ;
        END
        AntennaGateArea 0.169 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.095 -0.130 17.220 0.130 ;
        RECT  16.835 -0.130 17.095 0.955 ;
        RECT  16.050 -0.130 16.835 0.130 ;
        RECT  15.840 -0.130 16.050 0.990 ;
        RECT  15.105 -0.130 15.840 0.250 ;
        RECT  3.150 -0.130 15.105 0.130 ;
        RECT  2.890 -0.130 3.150 0.260 ;
        RECT  0.700 -0.130 2.890 0.130 ;
        RECT  0.200 -0.130 0.700 0.300 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.095 2.740 17.220 3.000 ;
        RECT  16.835 1.800 17.095 3.000 ;
        RECT  15.980 2.740 16.835 3.000 ;
        RECT  15.380 2.570 15.980 3.000 ;
        RECT  10.120 2.740 15.380 3.000 ;
        RECT  9.860 2.620 10.120 3.000 ;
        RECT  9.010 2.740 9.860 3.000 ;
        RECT  8.750 2.620 9.010 3.000 ;
        RECT  6.940 2.740 8.750 3.000 ;
        RECT  6.000 2.620 6.940 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.910 1.185 16.035 1.445 ;
        RECT  15.750 1.185 15.910 2.285 ;
        RECT  15.660 1.185 15.750 1.445 ;
        RECT  14.905 2.125 15.750 2.285 ;
        RECT  15.500 0.475 15.660 1.445 ;
        RECT  15.320 1.685 15.570 1.945 ;
        RECT  14.890 0.475 15.500 0.635 ;
        RECT  15.435 1.185 15.500 1.445 ;
        RECT  15.215 0.815 15.320 0.975 ;
        RECT  15.215 1.685 15.320 1.845 ;
        RECT  15.055 0.815 15.215 1.845 ;
        RECT  14.945 1.255 15.055 1.515 ;
        RECT  14.745 2.125 14.905 2.455 ;
        RECT  14.705 0.355 14.890 0.635 ;
        RECT  14.375 2.295 14.745 2.455 ;
        RECT  14.390 0.355 14.705 0.555 ;
        RECT  14.535 1.565 14.680 1.825 ;
        RECT  14.375 0.765 14.535 2.115 ;
        RECT  12.430 0.355 14.390 0.515 ;
        RECT  14.230 0.765 14.375 0.925 ;
        RECT  13.655 1.955 14.375 2.115 ;
        RECT  14.110 2.295 14.375 2.515 ;
        RECT  14.050 1.515 14.195 1.775 ;
        RECT  12.820 2.295 14.110 2.455 ;
        RECT  13.890 0.695 14.050 1.775 ;
        RECT  12.250 0.695 13.890 0.855 ;
        RECT  13.495 1.035 13.655 2.115 ;
        RECT  11.910 1.035 13.495 1.195 ;
        RECT  13.050 1.865 13.495 2.025 ;
        RECT  12.280 1.815 12.540 2.005 ;
        RECT  11.780 1.845 12.280 2.005 ;
        RECT  12.020 2.185 12.280 2.440 ;
        RECT  12.090 0.310 12.250 0.855 ;
        RECT  3.670 0.310 12.090 0.470 ;
        RECT  9.570 2.270 12.020 2.440 ;
        RECT  11.750 0.650 11.910 1.195 ;
        RECT  11.620 1.845 11.780 2.090 ;
        RECT  6.730 0.650 11.750 0.810 ;
        RECT  10.050 1.930 11.620 2.090 ;
        RECT  11.410 0.990 11.570 1.250 ;
        RECT  10.050 0.990 11.410 1.150 ;
        RECT  9.890 0.990 10.050 2.090 ;
        RECT  9.800 1.455 9.890 1.715 ;
        RECT  9.380 1.025 9.710 1.185 ;
        RECT  9.310 2.270 9.570 2.560 ;
        RECT  9.220 1.025 9.380 2.090 ;
        RECT  8.440 2.270 9.310 2.440 ;
        RECT  9.110 1.840 9.220 2.090 ;
        RECT  8.560 1.840 9.110 2.000 ;
        RECT  8.560 0.990 8.610 1.150 ;
        RECT  8.400 0.990 8.560 2.000 ;
        RECT  8.280 2.270 8.440 2.480 ;
        RECT  8.350 0.990 8.400 1.150 ;
        RECT  8.100 1.840 8.400 2.000 ;
        RECT  7.760 2.300 8.280 2.480 ;
        RECT  7.940 1.840 8.100 2.120 ;
        RECT  7.760 1.180 7.840 1.440 ;
        RECT  7.600 1.180 7.760 2.480 ;
        RECT  7.560 1.180 7.600 1.440 ;
        RECT  5.820 2.280 7.600 2.440 ;
        RECT  7.260 1.660 7.420 2.100 ;
        RECT  5.920 1.940 7.260 2.100 ;
        RECT  6.360 0.650 6.730 0.840 ;
        RECT  6.200 0.650 6.360 1.760 ;
        RECT  6.100 1.600 6.200 1.760 ;
        RECT  5.760 0.650 5.920 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.200 0.650 5.760 0.810 ;
        RECT  4.750 1.360 5.760 1.520 ;
        RECT  1.665 2.400 5.660 2.560 ;
        RECT  4.070 0.650 4.900 0.810 ;
        RECT  2.005 2.060 4.820 2.220 ;
        RECT  4.590 1.360 4.750 1.880 ;
        RECT  4.020 0.650 4.070 1.035 ;
        RECT  3.910 0.650 4.020 1.540 ;
        RECT  3.860 0.875 3.910 1.540 ;
        RECT  3.715 1.380 3.860 1.540 ;
        RECT  3.510 0.310 3.670 0.665 ;
        RECT  2.500 0.505 3.510 0.665 ;
        RECT  2.855 1.380 2.955 1.540 ;
        RECT  2.695 1.140 2.855 1.540 ;
        RECT  2.500 1.140 2.695 1.300 ;
        RECT  2.340 0.365 2.500 1.300 ;
        RECT  2.110 1.140 2.340 1.300 ;
        RECT  1.040 0.310 2.160 0.470 ;
        RECT  1.950 1.140 2.110 1.400 ;
        RECT  1.845 1.660 2.005 2.220 ;
        RECT  1.770 1.660 1.845 1.820 ;
        RECT  1.610 0.650 1.770 1.820 ;
        RECT  1.505 2.200 1.665 2.560 ;
        RECT  1.220 0.650 1.610 0.810 ;
        RECT  1.430 2.200 1.505 2.360 ;
        RECT  1.270 1.110 1.430 2.360 ;
        RECT  0.880 0.310 1.040 0.975 ;
        RECT  0.330 0.815 0.880 0.975 ;
        RECT  0.330 2.025 0.385 2.290 ;
        RECT  0.125 0.815 0.330 2.290 ;
    END
END SDFFSRHQX4MTH

MACRO SDFFSRHQX8MTH
    CLASS CORE ;
    FOREIGN SDFFSRHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.450 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 1.175 6.990 1.760 ;
        END
        AntennaGateArea 0.1807 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.270 2.060 5.480 2.220 ;
        RECT  5.020 1.700 5.270 2.220 ;
        END
        AntennaGateArea 0.0715 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.410 1.020 5.580 1.180 ;
        RECT  4.250 1.020 4.410 1.880 ;
        RECT  4.200 1.250 4.250 1.880 ;
        RECT  2.490 1.720 4.200 1.880 ;
        RECT  2.220 1.620 2.490 1.880 ;
        END
        AntennaGateArea 0.1287 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.055 1.385 13.315 1.635 ;
        RECT  11.010 1.440 13.055 1.635 ;
        RECT  10.540 1.330 11.010 1.635 ;
        END
        AntennaGateArea 0.2041 ;
    END RN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.500 0.400 17.760 2.285 ;
        RECT  16.650 1.290 17.500 1.580 ;
        RECT  16.390 0.400 16.650 2.285 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.080 0.875 3.640 1.180 ;
        END
        AntennaGateArea 0.13 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.470 1.235 0.760 1.830 ;
        END
        AntennaGateArea 0.169 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.310 -0.130 18.450 0.130 ;
        RECT  18.050 -0.130 18.310 1.025 ;
        RECT  17.205 -0.130 18.050 0.130 ;
        RECT  16.945 -0.130 17.205 1.025 ;
        RECT  16.100 -0.130 16.945 0.130 ;
        RECT  15.840 -0.130 16.100 1.025 ;
        RECT  3.150 -0.130 15.840 0.130 ;
        RECT  2.890 -0.130 3.150 0.260 ;
        RECT  0.700 -0.130 2.890 0.130 ;
        RECT  0.200 -0.130 0.700 0.300 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.310 2.740 18.450 3.000 ;
        RECT  18.050 1.785 18.310 3.000 ;
        RECT  17.200 2.740 18.050 3.000 ;
        RECT  16.940 1.780 17.200 3.000 ;
        RECT  15.945 2.740 16.940 3.000 ;
        RECT  15.345 2.570 15.945 3.000 ;
        RECT  11.150 2.740 15.345 3.000 ;
        RECT  10.890 2.620 11.150 3.000 ;
        RECT  10.120 2.740 10.890 3.000 ;
        RECT  9.860 2.620 10.120 3.000 ;
        RECT  9.010 2.740 9.860 3.000 ;
        RECT  8.750 2.620 9.010 3.000 ;
        RECT  7.385 2.740 8.750 3.000 ;
        RECT  6.785 2.620 7.385 3.000 ;
        RECT  6.600 2.740 6.785 3.000 ;
        RECT  6.000 2.620 6.600 3.000 ;
        RECT  0.815 2.740 6.000 3.000 ;
        RECT  0.215 2.570 0.815 3.000 ;
        RECT  0.000 2.740 0.215 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.910 1.205 16.035 1.465 ;
        RECT  15.750 1.205 15.910 2.285 ;
        RECT  15.660 1.205 15.750 1.465 ;
        RECT  14.950 2.125 15.750 2.285 ;
        RECT  15.500 0.355 15.660 1.465 ;
        RECT  15.320 1.685 15.570 1.945 ;
        RECT  12.430 0.355 15.500 0.515 ;
        RECT  15.435 1.205 15.500 1.465 ;
        RECT  15.215 0.815 15.320 0.975 ;
        RECT  15.215 1.685 15.320 1.845 ;
        RECT  15.055 0.815 15.215 1.845 ;
        RECT  14.945 1.155 15.055 1.415 ;
        RECT  14.790 2.125 14.950 2.405 ;
        RECT  13.080 2.245 14.790 2.405 ;
        RECT  14.400 1.465 14.680 1.725 ;
        RECT  14.400 0.725 14.640 0.885 ;
        RECT  14.240 0.725 14.400 2.065 ;
        RECT  13.655 1.905 14.240 2.065 ;
        RECT  13.900 0.695 14.060 1.725 ;
        RECT  12.250 0.695 13.900 0.855 ;
        RECT  13.495 1.035 13.655 2.065 ;
        RECT  11.910 1.035 13.495 1.195 ;
        RECT  13.050 1.865 13.495 2.025 ;
        RECT  12.820 2.245 13.080 2.455 ;
        RECT  12.280 1.815 12.540 2.005 ;
        RECT  10.660 1.845 12.280 2.005 ;
        RECT  12.020 2.185 12.280 2.440 ;
        RECT  12.090 0.310 12.250 0.855 ;
        RECT  3.670 0.310 12.090 0.470 ;
        RECT  9.570 2.270 12.020 2.440 ;
        RECT  11.750 0.650 11.910 1.195 ;
        RECT  6.730 0.650 11.750 0.810 ;
        RECT  11.410 0.990 11.570 1.250 ;
        RECT  10.050 0.990 11.410 1.150 ;
        RECT  10.400 1.845 10.660 2.090 ;
        RECT  10.050 1.845 10.400 2.005 ;
        RECT  9.890 0.990 10.050 2.005 ;
        RECT  9.800 1.455 9.890 1.715 ;
        RECT  9.380 1.025 9.710 1.185 ;
        RECT  9.310 2.270 9.570 2.560 ;
        RECT  9.220 1.025 9.380 2.090 ;
        RECT  8.440 2.270 9.310 2.440 ;
        RECT  9.110 1.840 9.220 2.090 ;
        RECT  8.350 1.840 9.110 2.000 ;
        RECT  8.350 0.990 8.610 1.150 ;
        RECT  8.280 2.270 8.440 2.490 ;
        RECT  8.190 0.990 8.350 2.000 ;
        RECT  7.760 2.300 8.280 2.490 ;
        RECT  8.100 1.840 8.190 2.000 ;
        RECT  7.940 1.840 8.100 2.120 ;
        RECT  7.760 1.180 7.840 1.440 ;
        RECT  7.600 1.180 7.760 2.490 ;
        RECT  7.555 1.180 7.600 1.440 ;
        RECT  5.820 2.280 7.600 2.440 ;
        RECT  7.260 1.695 7.420 2.100 ;
        RECT  5.920 1.940 7.260 2.100 ;
        RECT  6.360 0.650 6.730 0.840 ;
        RECT  6.200 0.650 6.360 1.760 ;
        RECT  6.100 1.600 6.200 1.760 ;
        RECT  5.760 0.650 5.920 2.100 ;
        RECT  5.660 2.280 5.820 2.560 ;
        RECT  5.210 0.650 5.760 0.810 ;
        RECT  4.750 1.360 5.760 1.520 ;
        RECT  1.665 2.400 5.660 2.560 ;
        RECT  4.070 0.650 4.900 0.810 ;
        RECT  2.005 2.060 4.840 2.220 ;
        RECT  4.590 1.360 4.750 1.880 ;
        RECT  4.020 0.650 4.070 1.035 ;
        RECT  3.910 0.650 4.020 1.540 ;
        RECT  3.860 0.875 3.910 1.540 ;
        RECT  3.715 1.380 3.860 1.540 ;
        RECT  3.510 0.310 3.670 0.665 ;
        RECT  2.500 0.505 3.510 0.665 ;
        RECT  2.855 1.380 2.955 1.540 ;
        RECT  2.695 1.135 2.855 1.540 ;
        RECT  2.500 1.135 2.695 1.295 ;
        RECT  2.340 0.365 2.500 1.295 ;
        RECT  2.110 1.135 2.340 1.295 ;
        RECT  1.040 0.310 2.160 0.470 ;
        RECT  1.950 1.135 2.110 1.400 ;
        RECT  1.845 1.860 2.005 2.220 ;
        RECT  1.770 1.860 1.845 2.020 ;
        RECT  1.610 0.650 1.770 2.020 ;
        RECT  1.505 2.200 1.665 2.560 ;
        RECT  1.220 0.650 1.610 0.810 ;
        RECT  1.100 2.200 1.505 2.360 ;
        RECT  1.270 1.110 1.430 1.370 ;
        RECT  1.100 1.210 1.270 1.370 ;
        RECT  0.940 1.210 1.100 2.360 ;
        RECT  0.880 0.310 1.040 0.790 ;
        RECT  0.385 0.630 0.880 0.790 ;
        RECT  0.285 0.630 0.385 1.025 ;
        RECT  0.285 2.030 0.385 2.290 ;
        RECT  0.125 0.630 0.285 2.290 ;
    END
END SDFFSRHQX8MTH

MACRO SDFFSRX1MTH
    CLASS CORE ;
    FOREIGN SDFFSRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.170 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.270 1.805 12.530 2.405 ;
        RECT  11.990 2.110 12.270 2.405 ;
        END
        AntennaGateArea 0.1118 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.480 1.975 2.100 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 1.155 1.200 1.540 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.820 1.330 6.500 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.495 0.640 14.655 2.045 ;
        RECT  13.845 0.640 14.495 0.800 ;
        RECT  14.250 1.885 14.495 2.045 ;
        RECT  13.790 1.885 14.250 2.400 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.835 0.755 15.070 2.120 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.545 1.110 1.965 1.270 ;
        RECT  1.385 1.110 1.545 2.100 ;
        RECT  1.285 1.700 1.385 2.100 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.400 1.110 5.640 1.580 ;
        RECT  5.355 1.190 5.400 1.450 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.985 -0.130 15.170 0.130 ;
        RECT  14.385 -0.130 14.985 0.345 ;
        RECT  13.150 -0.130 14.385 0.130 ;
        RECT  12.890 -0.130 13.150 0.345 ;
        RECT  6.020 -0.130 12.890 0.130 ;
        RECT  5.420 -0.130 6.020 0.250 ;
        RECT  4.710 -0.130 5.420 0.130 ;
        RECT  4.110 -0.130 4.710 0.250 ;
        RECT  1.855 -0.130 4.110 0.130 ;
        RECT  1.255 -0.130 1.855 0.250 ;
        RECT  0.955 -0.130 1.255 0.130 ;
        RECT  0.695 -0.130 0.955 0.250 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.475 2.740 15.170 3.000 ;
        RECT  14.215 2.580 14.475 3.000 ;
        RECT  13.440 2.740 14.215 3.000 ;
        RECT  13.280 1.905 13.440 3.000 ;
        RECT  4.045 2.740 13.280 3.000 ;
        RECT  3.885 2.245 4.045 3.000 ;
        RECT  1.745 2.740 3.885 3.000 ;
        RECT  1.485 2.620 1.745 3.000 ;
        RECT  0.335 2.740 1.485 3.000 ;
        RECT  0.175 1.760 0.335 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.155 1.315 14.315 1.625 ;
        RECT  13.635 1.465 14.155 1.625 ;
        RECT  13.475 0.605 13.635 1.625 ;
        RECT  13.320 0.605 13.475 0.765 ;
        RECT  12.870 1.465 13.475 1.625 ;
        RECT  13.030 0.960 13.290 1.255 ;
        RECT  10.270 1.095 13.030 1.255 ;
        RECT  12.710 1.465 12.870 1.945 ;
        RECT  11.220 1.465 12.710 1.625 ;
        RECT  12.400 0.310 12.560 0.760 ;
        RECT  10.715 0.310 12.400 0.470 ;
        RECT  9.930 0.755 11.920 0.915 ;
        RECT  11.590 2.015 11.690 2.175 ;
        RECT  11.430 2.015 11.590 2.560 ;
        RECT  7.920 2.400 11.430 2.560 ;
        RECT  10.610 1.595 10.950 1.855 ;
        RECT  10.115 0.310 10.715 0.575 ;
        RECT  10.450 1.595 10.610 2.220 ;
        RECT  8.800 2.060 10.450 2.220 ;
        RECT  10.110 1.095 10.270 1.880 ;
        RECT  9.100 0.310 10.115 0.470 ;
        RECT  9.760 1.720 10.110 1.880 ;
        RECT  9.770 0.755 9.930 1.540 ;
        RECT  9.230 1.380 9.770 1.540 ;
        RECT  9.430 0.655 9.590 1.200 ;
        RECT  8.180 1.040 9.430 1.200 ;
        RECT  9.110 1.380 9.230 1.570 ;
        RECT  8.950 1.380 9.110 1.760 ;
        RECT  8.840 0.310 9.100 0.860 ;
        RECT  7.535 1.600 8.950 1.760 ;
        RECT  8.640 1.955 8.800 2.220 ;
        RECT  7.480 1.955 8.640 2.115 ;
        RECT  8.060 1.040 8.180 1.420 ;
        RECT  7.900 0.310 8.060 1.420 ;
        RECT  7.660 2.295 7.920 2.560 ;
        RECT  6.360 0.310 7.900 0.470 ;
        RECT  7.375 0.650 7.535 1.760 ;
        RECT  7.320 1.955 7.480 2.220 ;
        RECT  4.385 2.400 7.480 2.560 ;
        RECT  6.700 0.650 7.375 0.810 ;
        RECT  4.725 2.060 7.320 2.220 ;
        RECT  6.965 0.990 7.150 1.880 ;
        RECT  6.890 0.990 6.965 1.150 ;
        RECT  6.000 1.720 6.965 1.880 ;
        RECT  6.540 0.650 6.700 0.930 ;
        RECT  5.175 0.770 6.540 0.930 ;
        RECT  6.200 0.310 6.360 0.590 ;
        RECT  4.105 0.430 6.200 0.590 ;
        RECT  5.175 1.720 5.285 1.880 ;
        RECT  5.015 0.770 5.175 1.880 ;
        RECT  4.785 1.110 5.015 1.270 ;
        RECT  4.445 0.770 4.835 0.930 ;
        RECT  4.625 1.110 4.785 1.370 ;
        RECT  4.565 1.565 4.725 2.220 ;
        RECT  4.445 1.565 4.565 1.725 ;
        RECT  4.285 0.770 4.445 1.725 ;
        RECT  4.225 1.905 4.385 2.560 ;
        RECT  3.625 1.565 4.285 1.725 ;
        RECT  3.375 1.905 4.225 2.065 ;
        RECT  3.945 0.430 4.105 1.100 ;
        RECT  3.465 0.785 3.625 1.725 ;
        RECT  2.995 1.545 3.465 1.725 ;
        RECT  3.215 1.905 3.375 2.175 ;
        RECT  3.095 0.635 3.255 1.365 ;
        RECT  2.655 2.015 3.215 2.175 ;
        RECT  2.655 1.205 3.095 1.365 ;
        RECT  2.835 1.545 2.995 1.835 ;
        RECT  2.315 0.770 2.735 0.975 ;
        RECT  2.495 1.205 2.655 2.175 ;
        RECT  2.315 2.355 2.635 2.515 ;
        RECT  2.275 0.360 2.535 0.590 ;
        RECT  2.155 0.770 2.315 2.515 ;
        RECT  0.525 0.430 2.275 0.590 ;
        RECT  0.970 0.770 2.155 0.930 ;
        RECT  0.895 2.280 2.155 2.440 ;
        RECT  0.705 0.770 0.970 0.960 ;
        RECT  0.675 1.735 0.955 1.895 ;
        RECT  0.635 2.280 0.895 2.465 ;
        RECT  0.525 1.370 0.675 1.895 ;
        RECT  0.515 0.430 0.525 1.895 ;
        RECT  0.365 0.430 0.515 1.530 ;
        RECT  0.125 0.430 0.365 0.590 ;
    END
END SDFFSRX1MTH

MACRO SDFFSRX2MTH
    CLASS CORE ;
    FOREIGN SDFFSRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.170 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.270 1.820 12.530 2.420 ;
        RECT  11.990 2.110 12.270 2.420 ;
        END
        AntennaGateArea 0.1352 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.480 1.975 2.100 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 1.155 1.200 1.540 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.820 1.330 6.500 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.975 1.685 14.295 1.950 ;
        RECT  13.785 0.765 13.975 1.950 ;
        END
        AntennaDiffArea 0.511 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.835 0.425 15.070 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.545 1.110 1.965 1.270 ;
        RECT  1.385 1.110 1.545 2.100 ;
        RECT  1.285 1.700 1.385 2.100 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.400 1.110 5.640 1.580 ;
        RECT  5.355 1.190 5.400 1.450 ;
        END
        AntennaGateArea 0.1183 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.535 -0.130 15.170 0.130 ;
        RECT  14.275 -0.130 14.535 0.955 ;
        RECT  6.020 -0.130 14.275 0.130 ;
        RECT  5.420 -0.130 6.020 0.250 ;
        RECT  5.035 -0.130 5.420 0.130 ;
        RECT  4.095 -0.130 5.035 0.250 ;
        RECT  1.855 -0.130 4.095 0.130 ;
        RECT  1.255 -0.130 1.855 0.250 ;
        RECT  0.955 -0.130 1.255 0.130 ;
        RECT  0.695 -0.130 0.955 0.250 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.505 2.740 15.170 3.000 ;
        RECT  14.245 2.470 14.505 3.000 ;
        RECT  13.455 2.740 14.245 3.000 ;
        RECT  12.855 2.470 13.455 3.000 ;
        RECT  4.045 2.740 12.855 3.000 ;
        RECT  3.885 2.245 4.045 3.000 ;
        RECT  1.745 2.740 3.885 3.000 ;
        RECT  1.485 2.620 1.745 3.000 ;
        RECT  0.335 2.740 1.485 3.000 ;
        RECT  0.175 1.760 0.335 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.495 1.245 14.655 2.290 ;
        RECT  13.580 2.130 14.495 2.290 ;
        RECT  13.420 0.355 13.580 2.290 ;
        RECT  13.320 0.355 13.420 0.515 ;
        RECT  12.870 1.825 13.420 1.985 ;
        RECT  13.080 1.095 13.240 1.465 ;
        RECT  10.270 1.095 13.080 1.255 ;
        RECT  12.710 1.465 12.870 1.985 ;
        RECT  11.220 1.465 12.710 1.625 ;
        RECT  12.400 0.310 12.560 0.785 ;
        RECT  10.715 0.310 12.400 0.470 ;
        RECT  9.930 0.755 11.925 0.915 ;
        RECT  11.590 2.015 11.690 2.175 ;
        RECT  11.430 2.015 11.590 2.560 ;
        RECT  7.920 2.400 11.430 2.560 ;
        RECT  10.610 1.595 10.950 1.855 ;
        RECT  10.115 0.310 10.715 0.575 ;
        RECT  10.450 1.595 10.610 2.220 ;
        RECT  8.800 2.060 10.450 2.220 ;
        RECT  10.110 1.095 10.270 1.880 ;
        RECT  9.100 0.310 10.115 0.470 ;
        RECT  9.760 1.720 10.110 1.880 ;
        RECT  9.770 0.755 9.930 1.540 ;
        RECT  9.240 1.380 9.770 1.540 ;
        RECT  9.430 0.655 9.590 1.200 ;
        RECT  8.180 1.040 9.430 1.200 ;
        RECT  9.120 1.380 9.240 1.615 ;
        RECT  8.960 1.380 9.120 1.760 ;
        RECT  8.930 0.310 9.100 0.830 ;
        RECT  7.535 1.600 8.960 1.760 ;
        RECT  8.840 0.670 8.930 0.830 ;
        RECT  8.640 1.955 8.800 2.220 ;
        RECT  7.480 1.955 8.640 2.115 ;
        RECT  8.060 1.040 8.180 1.420 ;
        RECT  7.900 0.310 8.060 1.420 ;
        RECT  7.660 2.295 7.920 2.560 ;
        RECT  6.360 0.310 7.900 0.470 ;
        RECT  7.375 0.650 7.535 1.760 ;
        RECT  7.320 1.955 7.480 2.220 ;
        RECT  4.385 2.400 7.480 2.560 ;
        RECT  6.700 0.650 7.375 0.810 ;
        RECT  4.725 2.060 7.320 2.220 ;
        RECT  6.955 0.990 7.150 1.880 ;
        RECT  6.890 0.990 6.955 1.150 ;
        RECT  6.000 1.720 6.955 1.880 ;
        RECT  6.540 0.650 6.700 0.930 ;
        RECT  5.175 0.770 6.540 0.930 ;
        RECT  6.200 0.310 6.360 0.590 ;
        RECT  4.105 0.430 6.200 0.590 ;
        RECT  5.175 1.720 5.285 1.880 ;
        RECT  5.015 0.770 5.175 1.880 ;
        RECT  4.785 1.110 5.015 1.270 ;
        RECT  4.445 0.770 4.835 0.930 ;
        RECT  4.625 1.110 4.785 1.370 ;
        RECT  4.565 1.565 4.725 2.220 ;
        RECT  4.445 1.565 4.565 1.725 ;
        RECT  4.285 0.770 4.445 1.725 ;
        RECT  4.225 1.905 4.385 2.560 ;
        RECT  3.625 1.565 4.285 1.725 ;
        RECT  3.375 1.905 4.225 2.065 ;
        RECT  3.945 0.430 4.105 1.100 ;
        RECT  3.465 0.785 3.625 1.725 ;
        RECT  2.995 1.545 3.465 1.725 ;
        RECT  3.215 1.905 3.375 2.175 ;
        RECT  3.095 0.635 3.255 1.365 ;
        RECT  3.205 2.015 3.215 2.175 ;
        RECT  2.945 2.015 3.205 2.275 ;
        RECT  2.655 1.205 3.095 1.365 ;
        RECT  2.835 1.545 2.995 1.835 ;
        RECT  2.655 2.015 2.945 2.175 ;
        RECT  2.315 0.770 2.735 0.945 ;
        RECT  2.495 1.205 2.655 2.175 ;
        RECT  2.315 2.355 2.635 2.515 ;
        RECT  2.275 0.360 2.535 0.590 ;
        RECT  2.155 0.770 2.315 2.515 ;
        RECT  0.525 0.430 2.275 0.590 ;
        RECT  0.965 0.770 2.155 0.930 ;
        RECT  0.895 2.280 2.155 2.440 ;
        RECT  0.705 0.770 0.965 0.960 ;
        RECT  0.675 1.735 0.955 1.895 ;
        RECT  0.635 2.280 0.895 2.465 ;
        RECT  0.525 1.370 0.675 1.895 ;
        RECT  0.515 0.430 0.525 1.895 ;
        RECT  0.365 0.430 0.515 1.530 ;
        RECT  0.125 0.430 0.365 0.590 ;
    END
END SDFFSRX2MTH

MACRO SDFFSRX4MTH
    CLASS CORE ;
    FOREIGN SDFFSRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.400 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.270 1.820 12.530 2.420 ;
        RECT  11.990 2.110 12.270 2.420 ;
        END
        AntennaGateArea 0.1521 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.480 1.975 2.100 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.870 1.155 1.200 1.540 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.820 1.330 6.500 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.535 0.390 14.695 1.990 ;
        RECT  14.370 1.700 14.535 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.790 1.290 15.890 1.580 ;
        RECT  15.555 0.425 15.790 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.545 1.110 1.965 1.270 ;
        RECT  1.385 1.110 1.545 2.100 ;
        RECT  1.285 1.700 1.385 2.100 ;
        END
        AntennaGateArea 0.0715 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  5.400 1.110 5.640 1.580 ;
        RECT  5.355 1.190 5.400 1.450 ;
        END
        AntennaGateArea 0.1443 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.275 -0.130 16.400 0.130 ;
        RECT  16.015 -0.130 16.275 0.955 ;
        RECT  15.255 -0.130 16.015 0.130 ;
        RECT  14.995 -0.130 15.255 0.955 ;
        RECT  14.205 -0.130 14.995 0.130 ;
        RECT  13.605 -0.130 14.205 0.300 ;
        RECT  13.160 -0.130 13.605 0.130 ;
        RECT  13.120 -0.130 13.160 0.345 ;
        RECT  12.860 -0.130 13.120 0.800 ;
        RECT  6.020 -0.130 12.860 0.130 ;
        RECT  5.420 -0.130 6.020 0.250 ;
        RECT  4.710 -0.130 5.420 0.130 ;
        RECT  4.110 -0.130 4.710 0.250 ;
        RECT  1.855 -0.130 4.110 0.130 ;
        RECT  1.255 -0.130 1.855 0.250 ;
        RECT  0.955 -0.130 1.255 0.130 ;
        RECT  0.695 -0.130 0.955 0.250 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.275 2.740 16.400 3.000 ;
        RECT  16.015 1.865 16.275 3.000 ;
        RECT  15.195 2.740 16.015 3.000 ;
        RECT  14.935 2.525 15.195 3.000 ;
        RECT  13.835 2.740 14.935 3.000 ;
        RECT  13.235 2.200 13.835 3.000 ;
        RECT  4.045 2.740 13.235 3.000 ;
        RECT  3.885 2.245 4.045 3.000 ;
        RECT  1.745 2.740 3.885 3.000 ;
        RECT  1.485 2.620 1.745 3.000 ;
        RECT  0.335 2.740 1.485 3.000 ;
        RECT  0.175 1.760 0.335 3.000 ;
        RECT  0.000 2.740 0.175 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.215 1.285 15.375 2.330 ;
        RECT  14.190 2.170 15.215 2.330 ;
        RECT  14.030 0.750 14.190 2.330 ;
        RECT  13.370 0.750 14.030 0.910 ;
        RECT  12.870 1.785 14.030 1.945 ;
        RECT  13.160 1.095 13.760 1.460 ;
        RECT  10.270 1.095 13.160 1.255 ;
        RECT  12.710 1.465 12.870 1.945 ;
        RECT  11.220 1.465 12.710 1.625 ;
        RECT  12.350 0.310 12.610 0.905 ;
        RECT  10.715 0.310 12.350 0.470 ;
        RECT  9.930 0.755 11.920 0.915 ;
        RECT  11.590 2.015 11.690 2.175 ;
        RECT  11.430 2.015 11.590 2.560 ;
        RECT  7.920 2.400 11.430 2.560 ;
        RECT  10.610 1.595 10.950 1.855 ;
        RECT  10.115 0.310 10.715 0.575 ;
        RECT  10.450 1.595 10.610 2.220 ;
        RECT  8.800 2.060 10.450 2.220 ;
        RECT  10.110 1.095 10.270 1.880 ;
        RECT  9.100 0.310 10.115 0.470 ;
        RECT  9.760 1.720 10.110 1.880 ;
        RECT  9.770 0.755 9.930 1.540 ;
        RECT  9.270 1.380 9.770 1.540 ;
        RECT  9.430 0.655 9.590 1.200 ;
        RECT  8.180 1.040 9.430 1.200 ;
        RECT  9.150 1.380 9.270 1.615 ;
        RECT  8.990 1.380 9.150 1.760 ;
        RECT  8.930 0.310 9.100 0.860 ;
        RECT  7.535 1.600 8.990 1.760 ;
        RECT  8.840 0.700 8.930 0.860 ;
        RECT  8.640 1.955 8.800 2.220 ;
        RECT  7.480 1.955 8.640 2.115 ;
        RECT  8.060 1.040 8.180 1.420 ;
        RECT  7.900 0.310 8.060 1.420 ;
        RECT  7.660 2.295 7.920 2.560 ;
        RECT  6.360 0.310 7.900 0.470 ;
        RECT  7.375 0.650 7.535 1.760 ;
        RECT  7.320 1.955 7.480 2.220 ;
        RECT  4.385 2.400 7.480 2.560 ;
        RECT  6.700 0.650 7.375 0.810 ;
        RECT  4.725 2.060 7.320 2.220 ;
        RECT  6.930 0.990 7.150 1.880 ;
        RECT  6.890 0.990 6.930 1.150 ;
        RECT  6.000 1.720 6.930 1.880 ;
        RECT  6.540 0.650 6.700 0.930 ;
        RECT  5.175 0.770 6.540 0.930 ;
        RECT  6.200 0.310 6.360 0.590 ;
        RECT  4.105 0.430 6.200 0.590 ;
        RECT  5.175 1.720 5.285 1.880 ;
        RECT  5.015 0.770 5.175 1.880 ;
        RECT  4.785 1.110 5.015 1.270 ;
        RECT  4.445 0.770 4.835 0.930 ;
        RECT  4.625 1.110 4.785 1.370 ;
        RECT  4.565 1.565 4.725 2.220 ;
        RECT  4.445 1.565 4.565 1.725 ;
        RECT  4.285 0.770 4.445 1.725 ;
        RECT  4.225 1.905 4.385 2.560 ;
        RECT  3.625 1.565 4.285 1.725 ;
        RECT  3.545 1.905 4.225 2.065 ;
        RECT  3.945 0.430 4.105 1.100 ;
        RECT  3.465 0.785 3.625 1.725 ;
        RECT  3.385 1.905 3.545 2.175 ;
        RECT  2.995 1.545 3.465 1.725 ;
        RECT  2.655 2.015 3.385 2.175 ;
        RECT  3.095 0.635 3.255 1.365 ;
        RECT  2.655 1.205 3.095 1.365 ;
        RECT  2.835 1.545 2.995 1.835 ;
        RECT  2.315 0.770 2.735 0.945 ;
        RECT  2.495 1.205 2.655 2.175 ;
        RECT  2.315 2.355 2.635 2.515 ;
        RECT  2.275 0.345 2.535 0.590 ;
        RECT  2.155 0.770 2.315 2.515 ;
        RECT  0.525 0.430 2.275 0.590 ;
        RECT  0.965 0.770 2.155 0.930 ;
        RECT  0.895 2.280 2.155 2.440 ;
        RECT  0.705 0.770 0.965 0.955 ;
        RECT  0.675 1.735 0.955 1.895 ;
        RECT  0.635 2.280 0.895 2.465 ;
        RECT  0.525 1.370 0.675 1.895 ;
        RECT  0.515 0.430 0.525 1.895 ;
        RECT  0.365 0.430 0.515 1.530 ;
        RECT  0.125 0.430 0.365 0.590 ;
    END
END SDFFSRX4MTH

MACRO SDFFSX1MTH
    CLASS CORE ;
    FOREIGN SDFFSX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.800 1.330 9.370 1.620 ;
        RECT  8.620 1.460 8.800 1.620 ;
        RECT  8.460 1.460 8.620 2.490 ;
        RECT  7.915 2.330 8.460 2.490 ;
        END
        AntennaGateArea 0.1118 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.240 1.580 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 1.110 0.360 1.740 ;
        RECT  0.100 1.290 0.130 1.580 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.350 0.815 10.560 1.990 ;
        RECT  10.120 0.815 10.350 1.075 ;
        RECT  10.115 1.725 10.350 1.990 ;
        END
        AntennaDiffArea 0.344 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 0.740 11.380 2.020 ;
        RECT  11.220 0.740 11.355 2.070 ;
        RECT  11.095 0.740 11.220 1.000 ;
        RECT  11.170 1.700 11.220 2.070 ;
        RECT  11.095 1.810 11.170 2.070 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.025 2.270 1.305 ;
        RECT  1.950 1.145 2.110 1.305 ;
        RECT  1.790 1.145 1.950 1.990 ;
        RECT  1.740 1.700 1.790 1.990 ;
        RECT  1.285 1.770 1.740 1.990 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.320 4.805 1.510 ;
        RECT  4.160 1.320 4.450 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.125 -0.130 11.480 0.130 ;
        RECT  10.525 -0.130 11.125 0.250 ;
        RECT  9.010 -0.130 10.525 0.130 ;
        RECT  8.750 -0.130 9.010 0.300 ;
        RECT  8.300 -0.130 8.750 0.130 ;
        RECT  7.700 -0.130 8.300 0.250 ;
        RECT  4.435 -0.130 7.700 0.130 ;
        RECT  4.175 -0.130 4.435 0.250 ;
        RECT  0.725 -0.130 4.175 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.075 2.740 11.480 3.000 ;
        RECT  9.235 2.570 10.075 3.000 ;
        RECT  7.720 2.740 9.235 3.000 ;
        RECT  6.780 2.620 7.720 3.000 ;
        RECT  1.745 2.740 6.780 3.000 ;
        RECT  1.485 2.620 1.745 3.000 ;
        RECT  0.385 2.740 1.485 3.000 ;
        RECT  0.125 2.230 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.900 1.190 11.040 1.450 ;
        RECT  10.740 0.435 10.900 2.330 ;
        RECT  10.010 0.435 10.740 0.595 ;
        RECT  9.865 2.170 10.740 2.330 ;
        RECT  9.710 1.265 10.150 1.525 ;
        RECT  9.750 0.355 10.010 0.595 ;
        RECT  9.605 1.960 9.865 2.330 ;
        RECT  9.550 0.990 9.710 1.525 ;
        RECT  8.960 2.170 9.605 2.330 ;
        RECT  8.280 0.990 9.550 1.150 ;
        RECT  8.510 0.640 9.040 0.800 ;
        RECT  8.800 2.170 8.960 2.450 ;
        RECT  8.350 0.475 8.510 0.800 ;
        RECT  7.520 0.475 8.350 0.635 ;
        RECT  8.170 0.990 8.280 2.150 ;
        RECT  8.120 0.815 8.170 2.150 ;
        RECT  7.940 0.815 8.120 1.150 ;
        RECT  7.650 1.990 8.120 2.150 ;
        RECT  7.600 0.865 7.760 1.790 ;
        RECT  7.490 1.990 7.650 2.440 ;
        RECT  7.180 0.865 7.600 1.025 ;
        RECT  7.310 1.630 7.600 1.790 ;
        RECT  7.360 0.310 7.520 0.635 ;
        RECT  6.690 2.280 7.490 2.440 ;
        RECT  6.840 1.210 7.420 1.450 ;
        RECT  6.055 0.310 7.360 0.470 ;
        RECT  7.150 1.630 7.310 2.100 ;
        RECT  7.020 0.650 7.180 1.025 ;
        RECT  7.050 1.940 7.150 2.100 ;
        RECT  6.400 0.650 7.020 0.810 ;
        RECT  6.580 0.990 6.840 1.450 ;
        RECT  6.530 1.890 6.690 2.440 ;
        RECT  6.290 1.290 6.580 1.450 ;
        RECT  6.240 0.650 6.400 1.110 ;
        RECT  6.130 1.290 6.290 2.560 ;
        RECT  5.545 0.950 6.240 1.110 ;
        RECT  5.970 2.140 6.130 2.560 ;
        RECT  5.795 0.310 6.055 0.665 ;
        RECT  2.710 2.400 5.970 2.560 ;
        RECT  5.790 1.520 5.950 1.880 ;
        RECT  4.810 1.720 5.790 1.880 ;
        RECT  5.320 0.405 5.545 1.110 ;
        RECT  5.285 0.405 5.320 1.540 ;
        RECT  5.060 0.950 5.285 1.540 ;
        RECT  4.340 0.950 5.060 1.110 ;
        RECT  3.290 2.060 5.030 2.220 ;
        RECT  4.745 0.340 5.005 0.590 ;
        RECT  4.550 1.690 4.810 1.880 ;
        RECT  3.885 0.430 4.745 0.590 ;
        RECT  3.885 1.720 4.550 1.880 ;
        RECT  4.180 0.950 4.340 1.135 ;
        RECT  4.065 0.975 4.180 1.135 ;
        RECT  3.725 0.310 3.885 1.880 ;
        RECT  3.225 0.310 3.725 0.470 ;
        RECT  3.470 1.590 3.725 1.850 ;
        RECT  3.290 0.675 3.545 0.935 ;
        RECT  3.130 0.675 3.290 2.220 ;
        RECT  2.950 0.310 2.975 0.570 ;
        RECT  2.790 0.310 2.950 2.220 ;
        RECT  1.320 0.310 2.790 0.470 ;
        RECT  2.525 2.060 2.790 2.220 ;
        RECT  2.450 0.685 2.610 1.645 ;
        RECT  2.365 2.060 2.525 2.440 ;
        RECT  1.610 0.685 2.450 0.845 ;
        RECT  2.330 1.485 2.450 1.645 ;
        RECT  0.925 2.280 2.365 2.440 ;
        RECT  2.165 1.485 2.330 1.785 ;
        RECT  1.450 0.685 1.610 1.025 ;
        RECT  0.830 0.865 1.450 1.025 ;
        RECT  1.060 0.310 1.320 0.525 ;
        RECT  0.635 2.215 0.925 2.440 ;
        RECT  0.815 0.865 0.830 1.915 ;
        RECT  0.670 0.765 0.815 1.915 ;
        RECT  0.620 0.765 0.670 1.025 ;
        RECT  0.570 1.755 0.670 1.915 ;
    END
END SDFFSX1MTH

MACRO SDFFSX2MTH
    CLASS CORE ;
    FOREIGN SDFFSX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.800 1.330 9.380 1.620 ;
        RECT  8.640 1.460 8.800 1.620 ;
        RECT  8.480 1.460 8.640 2.560 ;
        RECT  7.880 2.400 8.480 2.560 ;
        END
        AntennaGateArea 0.1352 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.320 1.290 1.580 1.540 ;
        RECT  0.925 1.330 1.320 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.130 1.110 0.360 1.740 ;
        RECT  0.100 1.290 0.130 1.580 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.620 0.815 10.680 0.975 ;
        RECT  10.350 0.815 10.620 1.990 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.735 1.700 11.790 1.990 ;
        RECT  11.475 0.400 11.735 2.390 ;
        END
        AntennaDiffArea 0.541 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.025 2.270 1.305 ;
        RECT  1.950 1.145 2.110 1.305 ;
        RECT  1.790 1.145 1.950 1.990 ;
        RECT  1.730 1.700 1.790 1.990 ;
        RECT  1.285 1.770 1.730 1.990 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.450 1.320 4.805 1.510 ;
        RECT  4.160 1.320 4.450 1.540 ;
        END
        AntennaGateArea 0.1183 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.220 -0.130 11.890 0.130 ;
        RECT  10.960 -0.130 11.220 0.250 ;
        RECT  10.080 -0.130 10.960 0.130 ;
        RECT  9.480 -0.130 10.080 0.250 ;
        RECT  4.430 -0.130 9.480 0.130 ;
        RECT  4.170 -0.130 4.430 0.250 ;
        RECT  0.725 -0.130 4.170 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.190 2.740 11.890 3.000 ;
        RECT  10.930 2.570 11.190 3.000 ;
        RECT  9.880 2.740 10.930 3.000 ;
        RECT  8.940 2.570 9.880 3.000 ;
        RECT  7.695 2.740 8.940 3.000 ;
        RECT  6.755 2.620 7.695 3.000 ;
        RECT  1.745 2.740 6.755 3.000 ;
        RECT  1.485 2.620 1.745 3.000 ;
        RECT  0.385 2.740 1.485 3.000 ;
        RECT  0.125 2.230 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.110 1.190 11.290 1.450 ;
        RECT  11.080 0.435 11.110 1.450 ;
        RECT  10.920 0.435 11.080 2.375 ;
        RECT  10.170 0.435 10.920 0.595 ;
        RECT  10.140 2.215 10.920 2.375 ;
        RECT  9.910 0.435 10.170 0.830 ;
        RECT  9.810 1.265 10.170 1.525 ;
        RECT  9.880 1.870 10.140 2.375 ;
        RECT  8.980 2.215 9.880 2.375 ;
        RECT  9.650 0.990 9.810 1.525 ;
        RECT  8.300 0.990 9.650 1.150 ;
        RECT  8.935 0.310 9.195 0.790 ;
        RECT  8.820 2.095 8.980 2.375 ;
        RECT  6.085 0.310 8.935 0.470 ;
        RECT  8.140 0.815 8.300 2.130 ;
        RECT  8.095 0.815 8.140 1.075 ;
        RECT  8.040 1.940 8.140 2.130 ;
        RECT  7.630 1.970 8.040 2.130 ;
        RECT  7.635 0.845 7.795 1.790 ;
        RECT  7.480 0.845 7.635 1.025 ;
        RECT  7.280 1.630 7.635 1.790 ;
        RECT  7.470 1.970 7.630 2.440 ;
        RECT  7.320 0.650 7.480 1.025 ;
        RECT  6.690 2.280 7.470 2.440 ;
        RECT  7.085 1.210 7.455 1.450 ;
        RECT  6.515 0.650 7.320 0.810 ;
        RECT  7.120 1.630 7.280 2.100 ;
        RECT  7.020 1.940 7.120 2.100 ;
        RECT  6.825 0.990 7.085 1.450 ;
        RECT  6.290 1.290 6.825 1.450 ;
        RECT  6.530 1.930 6.690 2.440 ;
        RECT  6.355 0.650 6.515 1.110 ;
        RECT  5.515 0.950 6.355 1.110 ;
        RECT  6.130 1.290 6.290 2.560 ;
        RECT  5.970 2.135 6.130 2.560 ;
        RECT  5.825 0.310 6.085 0.520 ;
        RECT  2.710 2.400 5.970 2.560 ;
        RECT  5.790 1.530 5.950 1.880 ;
        RECT  4.810 1.720 5.790 1.880 ;
        RECT  5.320 0.360 5.515 1.110 ;
        RECT  5.255 0.360 5.320 1.540 ;
        RECT  5.060 0.770 5.255 1.540 ;
        RECT  4.325 0.770 5.060 0.930 ;
        RECT  3.290 2.060 5.030 2.220 ;
        RECT  4.745 0.340 5.005 0.590 ;
        RECT  4.550 1.690 4.810 1.880 ;
        RECT  3.885 0.430 4.745 0.590 ;
        RECT  3.885 1.720 4.550 1.880 ;
        RECT  4.165 0.770 4.325 1.140 ;
        RECT  4.065 0.980 4.165 1.140 ;
        RECT  3.725 0.430 3.885 1.880 ;
        RECT  3.415 0.430 3.725 0.590 ;
        RECT  3.470 1.590 3.725 1.850 ;
        RECT  3.385 0.770 3.545 1.030 ;
        RECT  3.155 0.310 3.415 0.590 ;
        RECT  3.290 0.870 3.385 1.030 ;
        RECT  3.130 0.870 3.290 2.220 ;
        RECT  2.950 0.430 2.975 0.690 ;
        RECT  2.790 0.310 2.950 2.220 ;
        RECT  1.315 0.310 2.790 0.470 ;
        RECT  2.525 2.060 2.790 2.220 ;
        RECT  2.450 0.685 2.610 1.645 ;
        RECT  2.365 2.060 2.525 2.440 ;
        RECT  1.610 0.685 2.450 0.845 ;
        RECT  2.330 1.485 2.450 1.645 ;
        RECT  0.925 2.280 2.365 2.440 ;
        RECT  2.165 1.485 2.330 1.785 ;
        RECT  1.450 0.685 1.610 1.025 ;
        RECT  0.815 0.865 1.450 1.025 ;
        RECT  1.055 0.310 1.315 0.545 ;
        RECT  0.635 2.215 0.925 2.440 ;
        RECT  0.700 1.755 0.865 1.915 ;
        RECT  0.700 0.765 0.815 1.025 ;
        RECT  0.540 0.765 0.700 1.915 ;
    END
END SDFFSX2MTH

MACRO SDFFSX4MTH
    CLASS CORE ;
    FOREIGN SDFFSX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.080 1.330 9.370 1.800 ;
        RECT  8.275 1.330 9.080 1.490 ;
        RECT  8.115 1.330 8.275 1.765 ;
        RECT  7.830 1.605 8.115 1.765 ;
        RECT  7.670 1.605 7.830 1.885 ;
        END
        AntennaGateArea 0.2002 ;
    END SN
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.200 1.240 1.540 1.605 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.305 0.565 1.580 ;
        RECT  0.100 1.035 0.360 1.755 ;
        END
        AntennaGateArea 0.1131 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.795 0.395 10.970 1.170 ;
        RECT  10.625 0.395 10.795 1.955 ;
        END
        AntennaDiffArea 0.608 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.110 1.290 12.200 1.580 ;
        RECT  11.775 0.405 12.110 2.400 ;
        END
        AntennaDiffArea 0.614 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.045 2.025 1.305 ;
        RECT  1.740 1.045 1.950 2.105 ;
        RECT  1.330 1.845 1.740 2.105 ;
        END
        AntennaGateArea 0.0624 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.020 0.830 4.515 1.130 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.550 -0.130 12.710 0.130 ;
        RECT  12.290 -0.130 12.550 0.990 ;
        RECT  11.520 -0.130 12.290 0.130 ;
        RECT  11.215 -0.130 11.520 0.990 ;
        RECT  10.140 -0.130 11.215 0.130 ;
        RECT  9.640 -0.130 10.140 0.300 ;
        RECT  9.445 -0.130 9.640 0.130 ;
        RECT  9.185 -0.130 9.445 0.640 ;
        RECT  3.910 -0.130 9.185 0.130 ;
        RECT  3.650 -0.130 3.910 0.250 ;
        RECT  0.385 -0.130 3.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.470 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.550 2.740 12.710 3.000 ;
        RECT  12.290 1.825 12.550 3.000 ;
        RECT  11.515 2.740 12.290 3.000 ;
        RECT  11.315 1.805 11.515 3.000 ;
        RECT  11.180 2.570 11.315 3.000 ;
        RECT  10.290 2.740 11.180 3.000 ;
        RECT  10.030 2.480 10.290 3.000 ;
        RECT  9.055 2.740 10.030 3.000 ;
        RECT  8.795 2.570 9.055 3.000 ;
        RECT  8.270 2.740 8.795 3.000 ;
        RECT  7.670 2.570 8.270 3.000 ;
        RECT  5.570 2.740 7.670 3.000 ;
        RECT  5.370 2.570 5.570 3.000 ;
        RECT  0.385 2.740 5.370 3.000 ;
        RECT  0.125 2.410 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.380 1.170 11.540 1.625 ;
        RECT  11.135 1.365 11.380 1.625 ;
        RECT  10.975 1.365 11.135 2.295 ;
        RECT  10.445 2.135 10.975 2.295 ;
        RECT  10.285 0.650 10.445 2.295 ;
        RECT  10.020 0.650 10.285 0.810 ;
        RECT  9.625 2.135 10.285 2.295 ;
        RECT  9.765 1.170 10.105 1.430 ;
        RECT  9.760 0.545 10.020 0.810 ;
        RECT  9.605 0.990 9.765 1.430 ;
        RECT  9.365 2.135 9.625 2.430 ;
        RECT  7.860 0.990 9.605 1.150 ;
        RECT  8.845 2.135 9.365 2.295 ;
        RECT  8.770 0.525 8.870 0.785 ;
        RECT  8.685 1.845 8.845 2.295 ;
        RECT  8.610 0.310 8.770 0.785 ;
        RECT  8.585 1.845 8.685 2.005 ;
        RECT  5.500 0.310 8.610 0.470 ;
        RECT  7.490 2.065 8.165 2.225 ;
        RECT  7.720 0.750 7.860 1.150 ;
        RECT  7.560 0.750 7.720 1.395 ;
        RECT  7.490 1.235 7.560 1.395 ;
        RECT  7.330 1.235 7.490 2.560 ;
        RECT  6.635 2.400 7.330 2.560 ;
        RECT  7.150 0.740 7.300 1.000 ;
        RECT  6.990 0.650 7.150 2.220 ;
        RECT  5.990 0.650 6.990 0.810 ;
        RECT  6.885 2.060 6.990 2.220 ;
        RECT  6.720 0.990 6.780 1.150 ;
        RECT  6.620 0.990 6.720 1.530 ;
        RECT  6.375 2.300 6.635 2.560 ;
        RECT  6.460 0.990 6.620 2.120 ;
        RECT  6.075 1.960 6.460 2.120 ;
        RECT  5.980 1.180 6.240 1.780 ;
        RECT  5.915 1.960 6.075 2.390 ;
        RECT  5.780 0.650 5.990 0.960 ;
        RECT  5.575 1.400 5.980 1.560 ;
        RECT  5.190 2.230 5.915 2.390 ;
        RECT  4.940 0.800 5.780 0.960 ;
        RECT  5.415 1.400 5.575 1.880 ;
        RECT  5.240 0.310 5.500 0.620 ;
        RECT  4.640 1.720 5.415 1.880 ;
        RECT  5.030 2.230 5.190 2.560 ;
        RECT  4.940 1.280 5.150 1.540 ;
        RECT  2.885 2.400 5.030 2.560 ;
        RECT  4.855 0.410 4.940 1.540 ;
        RECT  4.780 0.410 4.855 1.470 ;
        RECT  3.160 2.060 4.850 2.220 ;
        RECT  3.675 1.310 4.780 1.470 ;
        RECT  4.360 1.685 4.640 1.880 ;
        RECT  3.480 0.460 4.480 0.620 ;
        RECT  3.445 1.685 4.360 1.845 ;
        RECT  3.445 0.310 3.480 0.620 ;
        RECT  3.285 0.310 3.445 1.845 ;
        RECT  3.220 0.310 3.285 0.470 ;
        RECT  3.245 1.570 3.285 1.845 ;
        RECT  3.060 2.030 3.160 2.220 ;
        RECT  3.060 0.655 3.105 0.915 ;
        RECT  2.900 0.655 3.060 2.220 ;
        RECT  2.545 0.365 2.705 2.495 ;
        RECT  0.635 0.365 2.545 0.525 ;
        RECT  2.330 2.205 2.545 2.495 ;
        RECT  2.205 0.705 2.365 1.795 ;
        RECT  0.910 2.335 2.330 2.495 ;
        RECT  0.910 0.705 2.205 0.865 ;
        RECT  2.180 1.535 2.205 1.795 ;
        RECT  0.750 0.705 0.910 1.985 ;
        RECT  0.650 2.275 0.910 2.535 ;
        RECT  0.650 0.705 0.750 1.115 ;
        RECT  0.650 1.815 0.750 1.985 ;
    END
END SDFFSX4MTH

MACRO SDFFTRX1MTH
    CLASS CORE ;
    FOREIGN SDFFTRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 1.330 2.415 1.740 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.755 1.840 2.975 2.080 ;
        RECT  2.595 0.990 2.755 2.080 ;
        RECT  2.265 0.990 2.595 1.150 ;
        RECT  1.675 1.920 2.595 2.080 ;
        RECT  1.330 1.660 1.675 2.080 ;
        RECT  0.515 1.660 1.330 1.820 ;
        END
        AntennaGateArea 0.1456 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 0.880 3.590 1.170 ;
        RECT  3.275 0.310 3.435 1.170 ;
        RECT  1.415 0.310 3.275 0.470 ;
        RECT  1.255 0.310 1.415 1.030 ;
        RECT  0.905 0.870 1.255 1.030 ;
        END
        AntennaGateArea 0.0611 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.935 1.290 10.150 1.580 ;
        RECT  9.775 0.805 9.935 2.090 ;
        RECT  9.665 1.830 9.775 2.090 ;
        END
        AntennaDiffArea 0.342 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.810 0.735 10.970 2.115 ;
        RECT  10.760 0.735 10.810 1.170 ;
        RECT  10.685 1.855 10.810 2.115 ;
        RECT  10.685 0.735 10.760 0.995 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 2.400 1.195 2.560 ;
        RECT  0.935 2.110 1.150 2.560 ;
        RECT  0.730 2.110 0.935 2.400 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 0.880 4.410 1.320 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.820 -0.130 11.070 0.130 ;
        RECT  9.880 -0.130 10.820 0.250 ;
        RECT  9.030 -0.130 9.880 0.130 ;
        RECT  8.770 -0.130 9.030 0.250 ;
        RECT  7.170 -0.130 8.770 0.130 ;
        RECT  6.910 -0.130 7.170 0.730 ;
        RECT  4.570 -0.130 6.910 0.130 ;
        RECT  3.630 -0.130 4.570 0.250 ;
        RECT  0.955 -0.130 3.630 0.130 ;
        RECT  0.695 -0.130 0.955 0.660 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.435 2.740 11.070 3.000 ;
        RECT  10.175 1.825 10.435 3.000 ;
        RECT  9.345 2.740 10.175 3.000 ;
        RECT  8.405 2.620 9.345 3.000 ;
        RECT  6.620 2.740 8.405 3.000 ;
        RECT  6.460 2.050 6.620 3.000 ;
        RECT  4.245 2.740 6.460 3.000 ;
        RECT  3.985 2.620 4.245 3.000 ;
        RECT  2.765 2.740 3.985 3.000 ;
        RECT  2.505 2.620 2.765 3.000 ;
        RECT  0.755 2.740 2.505 3.000 ;
        RECT  0.155 2.620 0.755 3.000 ;
        RECT  0.000 2.740 0.155 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.505 1.315 10.615 1.575 ;
        RECT  10.345 0.465 10.505 1.575 ;
        RECT  9.610 0.465 10.345 0.625 ;
        RECT  9.580 0.355 9.610 0.625 ;
        RECT  9.420 0.355 9.580 1.485 ;
        RECT  9.350 0.355 9.420 0.515 ;
        RECT  9.365 1.325 9.420 1.485 ;
        RECT  9.205 1.325 9.365 2.235 ;
        RECT  9.070 0.765 9.230 1.145 ;
        RECT  8.625 1.635 9.205 1.795 ;
        RECT  8.230 0.765 9.070 0.925 ;
        RECT  8.465 1.465 8.625 1.795 ;
        RECT  8.070 0.495 8.230 2.115 ;
        RECT  7.050 2.400 8.190 2.560 ;
        RECT  7.730 1.955 8.070 2.115 ;
        RECT  7.520 0.655 7.680 1.080 ;
        RECT  7.430 0.920 7.520 1.080 ;
        RECT  7.270 0.920 7.430 2.065 ;
        RECT  6.910 0.920 7.270 1.080 ;
        RECT  6.890 1.360 7.050 2.560 ;
        RECT  6.750 0.920 6.910 1.180 ;
        RECT  6.570 1.360 6.890 1.520 ;
        RECT  6.230 1.700 6.710 1.860 ;
        RECT  6.410 0.325 6.570 1.520 ;
        RECT  5.090 0.325 6.410 0.485 ;
        RECT  6.070 0.685 6.230 1.860 ;
        RECT  5.850 1.700 6.070 1.860 ;
        RECT  5.690 1.700 5.850 2.340 ;
        RECT  5.460 0.705 5.710 0.865 ;
        RECT  5.450 2.180 5.690 2.340 ;
        RECT  5.300 0.705 5.460 2.000 ;
        RECT  5.090 1.840 5.300 2.000 ;
        RECT  4.930 0.325 5.090 1.660 ;
        RECT  4.930 1.840 5.090 2.420 ;
        RECT  4.595 1.500 4.930 1.660 ;
        RECT  3.655 2.260 4.930 2.420 ;
        RECT  4.590 0.480 4.750 1.180 ;
        RECT  4.435 1.500 4.595 1.860 ;
        RECT  3.930 0.480 4.590 0.640 ;
        RECT  3.770 0.480 3.930 1.795 ;
        RECT  3.655 1.635 3.770 1.795 ;
        RECT  3.495 1.635 3.655 1.895 ;
        RECT  3.395 2.260 3.655 2.475 ;
        RECT  3.315 2.260 3.395 2.420 ;
        RECT  3.155 1.415 3.315 2.420 ;
        RECT  3.095 1.415 3.155 1.575 ;
        RECT  1.875 2.260 3.155 2.420 ;
        RECT  2.935 0.650 3.095 1.575 ;
        RECT  1.895 0.650 2.935 0.810 ;
        RECT  1.745 1.100 1.905 1.480 ;
        RECT  1.615 2.260 1.875 2.475 ;
        RECT  0.335 1.320 1.745 1.480 ;
        RECT  0.175 0.570 0.335 2.240 ;
    END
END SDFFTRX1MTH

MACRO SDFFTRX2MTH
    CLASS CORE ;
    FOREIGN SDFFTRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.415 1.755 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.755 1.940 2.975 2.100 ;
        RECT  2.595 0.990 2.755 2.100 ;
        RECT  2.265 0.990 2.595 1.150 ;
        RECT  1.675 1.940 2.595 2.100 ;
        RECT  1.330 1.660 1.675 2.100 ;
        RECT  0.515 1.660 1.330 1.820 ;
        END
        AntennaGateArea 0.1456 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 0.880 3.590 1.170 ;
        RECT  3.275 0.310 3.435 1.170 ;
        RECT  1.415 0.310 3.275 0.470 ;
        RECT  1.255 0.310 1.415 1.030 ;
        RECT  0.905 0.870 1.255 1.030 ;
        END
        AntennaGateArea 0.0611 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.360 1.290 10.560 1.580 ;
        RECT  10.200 0.765 10.360 1.945 ;
        END
        AntennaDiffArea 0.497 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 0.420 11.380 1.170 ;
        RECT  11.195 0.420 11.355 2.425 ;
        RECT  11.170 0.420 11.195 1.170 ;
        RECT  11.095 1.825 11.195 2.425 ;
        RECT  11.095 0.420 11.170 1.020 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.150 2.400 1.195 2.560 ;
        RECT  0.935 2.110 1.150 2.560 ;
        RECT  0.730 2.110 0.935 2.400 ;
        END
        AntennaGateArea 0.0702 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 0.880 4.410 1.320 ;
        END
        AntennaGateArea 0.0975 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.435 -0.130 11.480 0.130 ;
        RECT  8.835 -0.130 9.435 0.250 ;
        RECT  7.170 -0.130 8.835 0.130 ;
        RECT  6.910 -0.130 7.170 0.575 ;
        RECT  4.570 -0.130 6.910 0.130 ;
        RECT  3.630 -0.130 4.570 0.250 ;
        RECT  0.955 -0.130 3.630 0.130 ;
        RECT  0.695 -0.130 0.955 0.660 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.390 2.740 11.480 3.000 ;
        RECT  8.790 2.620 9.390 3.000 ;
        RECT  7.630 2.740 8.790 3.000 ;
        RECT  7.470 2.245 7.630 3.000 ;
        RECT  6.550 2.740 7.470 3.000 ;
        RECT  6.390 2.050 6.550 3.000 ;
        RECT  4.245 2.740 6.390 3.000 ;
        RECT  3.985 2.620 4.245 3.000 ;
        RECT  2.765 2.740 3.985 3.000 ;
        RECT  2.505 2.620 2.765 3.000 ;
        RECT  0.755 2.740 2.505 3.000 ;
        RECT  0.155 2.620 0.755 3.000 ;
        RECT  0.000 2.740 0.155 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.900 1.305 11.010 1.565 ;
        RECT  10.740 0.355 10.900 1.565 ;
        RECT  9.990 0.355 10.740 0.515 ;
        RECT  9.830 0.355 9.990 1.525 ;
        RECT  9.480 2.245 9.970 2.405 ;
        RECT  9.640 0.525 9.830 0.685 ;
        RECT  9.480 1.365 9.830 1.525 ;
        RECT  9.490 0.885 9.650 1.145 ;
        RECT  9.140 0.985 9.490 1.145 ;
        RECT  9.320 1.365 9.480 2.405 ;
        RECT  8.980 0.985 9.140 2.300 ;
        RECT  8.530 0.985 8.980 1.145 ;
        RECT  8.330 2.140 8.980 2.300 ;
        RECT  8.640 1.365 8.800 1.695 ;
        RECT  8.190 1.365 8.640 1.525 ;
        RECT  8.370 0.465 8.530 1.145 ;
        RECT  8.030 0.355 8.190 1.525 ;
        RECT  7.850 1.785 8.080 1.945 ;
        RECT  7.510 0.355 8.030 0.515 ;
        RECT  7.690 0.765 7.850 1.945 ;
        RECT  7.090 1.095 7.690 1.255 ;
        RECT  7.350 0.355 7.510 0.915 ;
        RECT  6.570 0.755 7.350 0.915 ;
        RECT  6.930 1.095 7.090 2.155 ;
        RECT  6.700 1.095 6.930 1.255 ;
        RECT  6.230 1.575 6.750 1.735 ;
        RECT  6.410 0.325 6.570 0.915 ;
        RECT  5.090 0.325 6.410 0.485 ;
        RECT  6.070 0.685 6.230 1.735 ;
        RECT  5.850 1.575 6.070 1.735 ;
        RECT  5.690 1.575 5.850 2.340 ;
        RECT  5.460 0.705 5.710 0.865 ;
        RECT  5.450 2.180 5.690 2.340 ;
        RECT  5.300 0.705 5.460 2.000 ;
        RECT  5.090 1.840 5.300 2.000 ;
        RECT  4.930 0.325 5.090 1.660 ;
        RECT  4.930 1.840 5.090 2.440 ;
        RECT  4.595 1.500 4.930 1.660 ;
        RECT  3.655 2.280 4.930 2.440 ;
        RECT  4.590 0.540 4.750 1.180 ;
        RECT  4.435 1.500 4.595 1.860 ;
        RECT  3.930 0.540 4.590 0.700 ;
        RECT  3.770 0.540 3.930 1.795 ;
        RECT  3.655 1.635 3.770 1.795 ;
        RECT  3.495 1.635 3.655 1.895 ;
        RECT  3.395 2.280 3.655 2.475 ;
        RECT  3.315 2.280 3.395 2.440 ;
        RECT  3.155 1.525 3.315 2.440 ;
        RECT  3.095 1.525 3.155 1.685 ;
        RECT  1.875 2.280 3.155 2.440 ;
        RECT  2.935 0.650 3.095 1.685 ;
        RECT  1.895 0.650 2.935 0.810 ;
        RECT  1.745 1.100 1.905 1.480 ;
        RECT  1.615 2.280 1.875 2.475 ;
        RECT  0.335 1.320 1.745 1.480 ;
        RECT  0.175 0.570 0.335 2.240 ;
    END
END SDFFTRX2MTH

MACRO SDFFTRX4MTH
    CLASS CORE ;
    FOREIGN SDFFTRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.330 2.415 1.755 ;
        END
        AntennaGateArea 0.065 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.755 1.940 2.975 2.100 ;
        RECT  2.595 0.990 2.755 2.100 ;
        RECT  2.265 0.990 2.595 1.150 ;
        RECT  1.540 1.940 2.595 2.100 ;
        RECT  1.480 1.645 1.540 2.100 ;
        RECT  1.320 1.645 1.480 2.410 ;
        RECT  0.325 2.250 1.320 2.410 ;
        END
        AntennaGateArea 0.1885 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.435 0.880 3.590 1.170 ;
        RECT  3.275 0.310 3.435 1.170 ;
        RECT  1.415 0.310 3.275 0.470 ;
        RECT  1.255 0.310 1.415 1.060 ;
        RECT  0.905 0.900 1.255 1.060 ;
        END
        AntennaGateArea 0.0897 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.375 0.815 12.635 2.415 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.715 1.290 13.840 1.580 ;
        RECT  13.455 0.420 13.715 2.425 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.685 1.580 1.130 1.990 ;
        END
        AntennaGateArea 0.1248 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.110 0.880 4.410 1.320 ;
        END
        AntennaGateArea 0.1105 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 -0.130 14.350 0.130 ;
        RECT  13.965 -0.130 14.225 1.020 ;
        RECT  13.175 -0.130 13.965 0.130 ;
        RECT  12.915 -0.130 13.175 0.250 ;
        RECT  12.095 -0.130 12.915 0.130 ;
        RECT  11.835 -0.130 12.095 0.250 ;
        RECT  11.080 -0.130 11.835 0.130 ;
        RECT  10.480 -0.130 11.080 0.250 ;
        RECT  8.530 -0.130 10.480 0.130 ;
        RECT  8.370 -0.130 8.530 0.975 ;
        RECT  7.170 -0.130 8.370 0.130 ;
        RECT  6.910 -0.130 7.170 0.575 ;
        RECT  4.570 -0.130 6.910 0.130 ;
        RECT  3.630 -0.130 4.570 0.250 ;
        RECT  0.955 -0.130 3.630 0.130 ;
        RECT  0.695 -0.130 0.955 0.635 ;
        RECT  0.000 -0.130 0.695 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 2.740 14.350 3.000 ;
        RECT  13.965 1.825 14.225 3.000 ;
        RECT  13.175 2.740 13.965 3.000 ;
        RECT  12.915 1.825 13.175 3.000 ;
        RECT  12.125 2.740 12.915 3.000 ;
        RECT  11.865 1.825 12.125 3.000 ;
        RECT  11.105 2.740 11.865 3.000 ;
        RECT  10.845 1.845 11.105 3.000 ;
        RECT  10.475 2.325 10.845 3.000 ;
        RECT  8.590 2.740 10.475 3.000 ;
        RECT  8.430 1.955 8.590 3.000 ;
        RECT  7.570 2.740 8.430 3.000 ;
        RECT  7.410 1.920 7.570 3.000 ;
        RECT  6.550 2.740 7.410 3.000 ;
        RECT  6.390 1.955 6.550 3.000 ;
        RECT  4.245 2.740 6.390 3.000 ;
        RECT  3.985 2.620 4.245 3.000 ;
        RECT  2.765 2.740 3.985 3.000 ;
        RECT  2.505 2.620 2.765 3.000 ;
        RECT  0.865 2.740 2.505 3.000 ;
        RECT  0.265 2.620 0.865 3.000 ;
        RECT  0.000 2.740 0.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.115 0.475 13.275 1.485 ;
        RECT  11.975 0.475 13.115 0.635 ;
        RECT  11.815 0.475 11.975 0.965 ;
        RECT  11.565 0.805 11.815 0.965 ;
        RECT  11.565 1.935 11.615 2.195 ;
        RECT  11.405 0.805 11.565 2.195 ;
        RECT  11.240 0.395 11.500 0.590 ;
        RECT  10.970 1.135 11.405 1.295 ;
        RECT  11.355 1.935 11.405 2.195 ;
        RECT  10.630 0.430 11.240 0.590 ;
        RECT  10.810 1.135 10.970 1.395 ;
        RECT  10.470 0.430 10.630 2.055 ;
        RECT  10.030 0.800 10.470 0.960 ;
        RECT  10.160 1.895 10.470 2.055 ;
        RECT  10.130 1.225 10.290 1.705 ;
        RECT  10.000 1.895 10.160 2.505 ;
        RECT  9.550 1.225 10.130 1.385 ;
        RECT  9.770 0.700 10.030 0.960 ;
        RECT  9.150 2.345 10.000 2.505 ;
        RECT  9.450 1.565 9.610 2.125 ;
        RECT  9.390 0.395 9.550 1.385 ;
        RECT  9.210 1.565 9.450 1.725 ;
        RECT  8.870 0.395 9.390 0.555 ;
        RECT  9.050 0.785 9.210 1.725 ;
        RECT  8.890 1.945 9.150 2.505 ;
        RECT  8.080 1.565 9.050 1.725 ;
        RECT  8.710 0.395 8.870 1.385 ;
        RECT  8.190 1.225 8.710 1.385 ;
        RECT  8.030 0.545 8.190 1.385 ;
        RECT  7.920 1.565 8.080 2.180 ;
        RECT  7.510 0.545 8.030 0.705 ;
        RECT  7.850 1.565 7.920 1.725 ;
        RECT  7.690 0.895 7.850 1.725 ;
        RECT  7.060 1.095 7.690 1.255 ;
        RECT  7.350 0.545 7.510 0.915 ;
        RECT  6.540 0.755 7.350 0.915 ;
        RECT  6.900 1.095 7.060 2.180 ;
        RECT  6.700 1.095 6.900 1.255 ;
        RECT  6.200 1.575 6.710 1.735 ;
        RECT  6.380 0.325 6.540 0.915 ;
        RECT  5.170 0.325 6.380 0.485 ;
        RECT  6.040 0.685 6.200 1.735 ;
        RECT  5.850 1.575 6.040 1.735 ;
        RECT  5.690 1.575 5.850 2.340 ;
        RECT  5.510 0.705 5.740 0.865 ;
        RECT  5.450 2.180 5.690 2.340 ;
        RECT  5.350 0.705 5.510 2.000 ;
        RECT  5.120 1.840 5.350 2.000 ;
        RECT  5.010 0.325 5.170 1.660 ;
        RECT  4.960 1.840 5.120 2.440 ;
        RECT  4.930 0.550 5.010 0.810 ;
        RECT  4.610 1.500 5.010 1.660 ;
        RECT  3.655 2.280 4.960 2.440 ;
        RECT  4.590 0.540 4.750 1.180 ;
        RECT  4.450 1.500 4.610 1.860 ;
        RECT  3.930 0.540 4.590 0.700 ;
        RECT  3.770 0.540 3.930 1.795 ;
        RECT  3.655 1.635 3.770 1.795 ;
        RECT  3.495 1.635 3.655 1.895 ;
        RECT  3.395 2.280 3.655 2.480 ;
        RECT  3.315 2.280 3.395 2.440 ;
        RECT  3.155 1.525 3.315 2.440 ;
        RECT  3.095 1.525 3.155 1.685 ;
        RECT  1.825 2.280 3.155 2.440 ;
        RECT  2.935 0.650 3.095 1.685 ;
        RECT  1.895 0.650 2.935 0.810 ;
        RECT  1.745 1.140 1.905 1.400 ;
        RECT  1.665 2.280 1.825 2.540 ;
        RECT  0.335 1.240 1.745 1.400 ;
        RECT  0.335 1.880 0.385 2.040 ;
        RECT  0.175 0.600 0.335 2.040 ;
        RECT  0.125 1.880 0.175 2.040 ;
    END
END SDFFTRX4MTH

MACRO SDFFX1MTH
    CLASS CORE ;
    FOREIGN SDFFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.250 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.615 1.575 2.135 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 1.690 1.950 1.950 ;
        RECT  1.760 1.275 1.920 1.950 ;
        RECT  1.130 1.275 1.760 1.435 ;
        RECT  0.555 1.275 1.130 1.580 ;
        END
        AntennaGateArea 0.1261 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.665 0.875 8.825 1.135 ;
        RECT  8.510 2.355 8.760 2.515 ;
        RECT  8.225 0.975 8.665 1.135 ;
        RECT  8.300 2.110 8.510 2.515 ;
        RECT  8.225 2.110 8.300 2.270 ;
        RECT  8.065 0.975 8.225 2.270 ;
        END
        AntennaDiffArea 0.369 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.125 1.290 10.150 1.580 ;
        RECT  10.100 0.525 10.125 1.580 ;
        RECT  10.100 1.935 10.125 2.195 ;
        RECT  9.940 0.525 10.100 2.195 ;
        RECT  9.535 0.525 9.940 0.685 ;
        RECT  9.865 1.935 9.940 2.195 ;
        RECT  9.375 0.365 9.535 0.685 ;
        END
        AntennaDiffArea 0.316 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.100 2.360 1.580 ;
        END
        AntennaGateArea 0.0728 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.715 4.560 2.065 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.125 -0.130 10.250 0.130 ;
        RECT  9.865 -0.130 10.125 0.315 ;
        RECT  8.810 -0.130 9.865 0.130 ;
        RECT  7.870 -0.130 8.810 0.350 ;
        RECT  6.605 -0.130 7.870 0.130 ;
        RECT  6.345 -0.130 6.605 0.350 ;
        RECT  0.385 -0.130 6.345 0.130 ;
        RECT  0.125 -0.130 0.385 0.365 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.585 2.740 10.250 3.000 ;
        RECT  9.325 2.275 9.585 3.000 ;
        RECT  4.150 2.740 9.325 3.000 ;
        RECT  3.890 2.620 4.150 3.000 ;
        RECT  0.000 2.740 3.890 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.345 0.875 9.505 1.930 ;
        RECT  9.125 1.770 9.345 1.930 ;
        RECT  9.005 0.535 9.165 1.590 ;
        RECT  8.865 1.770 9.125 2.055 ;
        RECT  7.885 0.535 9.005 0.695 ;
        RECT  8.565 1.770 8.865 1.930 ;
        RECT  8.405 1.540 8.565 1.930 ;
        RECT  7.725 0.535 7.885 2.435 ;
        RECT  7.225 0.685 7.725 0.845 ;
        RECT  7.170 2.275 7.725 2.435 ;
        RECT  7.385 1.025 7.545 2.025 ;
        RECT  6.975 1.865 7.385 2.025 ;
        RECT  6.950 0.310 7.285 0.470 ;
        RECT  6.815 1.865 6.975 2.545 ;
        RECT  6.790 0.310 6.950 1.155 ;
        RECT  4.690 2.385 6.815 2.545 ;
        RECT  6.630 1.335 6.805 1.495 ;
        RECT  6.125 0.995 6.790 1.155 ;
        RECT  6.470 1.335 6.630 2.205 ;
        RECT  5.580 2.045 6.470 2.205 ;
        RECT  6.040 1.705 6.140 1.865 ;
        RECT  6.040 0.325 6.125 1.155 ;
        RECT  5.880 0.325 6.040 1.865 ;
        RECT  3.165 0.325 5.880 0.485 ;
        RECT  5.420 0.735 5.580 2.205 ;
        RECT  5.415 1.375 5.420 2.205 ;
        RECT  3.780 1.375 5.415 1.535 ;
        RECT  3.310 1.035 5.240 1.195 ;
        RECT  4.530 2.280 4.690 2.545 ;
        RECT  2.970 0.665 4.545 0.825 ;
        RECT  3.655 2.280 4.530 2.440 ;
        RECT  3.495 2.280 3.655 2.560 ;
        RECT  3.300 2.345 3.495 2.560 ;
        RECT  3.150 1.035 3.310 2.165 ;
        RECT  2.970 2.345 3.300 2.505 ;
        RECT  2.950 1.035 3.150 1.195 ;
        RECT  2.810 0.665 2.970 0.855 ;
        RECT  2.810 1.545 2.970 2.505 ;
        RECT  2.770 0.695 2.810 0.855 ;
        RECT  2.770 1.545 2.810 1.705 ;
        RECT  2.610 0.695 2.770 1.705 ;
        RECT  0.675 0.355 2.630 0.515 ;
        RECT  2.470 1.905 2.630 2.545 ;
        RECT  0.945 2.385 2.470 2.545 ;
        RECT  0.930 0.695 1.950 0.855 ;
        RECT  0.785 2.245 0.945 2.545 ;
        RECT  0.770 0.695 0.930 1.075 ;
        RECT  0.505 1.785 0.830 1.945 ;
        RECT  0.670 0.815 0.770 1.075 ;
        RECT  0.375 0.915 0.670 1.075 ;
        RECT  0.505 2.400 0.605 2.560 ;
        RECT  0.375 1.785 0.505 2.560 ;
        RECT  0.345 0.915 0.375 2.560 ;
        RECT  0.215 0.915 0.345 1.945 ;
    END
END SDFFX1MTH

MACRO SDFFX2MTH
    CLASS CORE ;
    FOREIGN SDFFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.615 1.575 2.135 ;
        RECT  1.125 1.760 1.310 2.135 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 1.925 1.950 2.185 ;
        RECT  1.760 1.275 1.920 2.185 ;
        RECT  1.130 1.275 1.760 1.435 ;
        RECT  0.685 1.275 1.130 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 1.290 10.560 1.580 ;
        RECT  10.275 0.400 10.535 2.355 ;
        END
        AntennaDiffArea 0.524 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.625 1.290 9.740 1.580 ;
        RECT  9.595 1.290 9.625 1.945 ;
        RECT  9.335 0.765 9.595 1.945 ;
        END
        AntennaDiffArea 0.42 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.100 2.360 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.160 1.715 4.560 2.065 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.995 -0.130 10.660 0.130 ;
        RECT  9.735 -0.130 9.995 0.515 ;
        RECT  8.970 -0.130 9.735 0.130 ;
        RECT  8.370 -0.130 8.970 0.250 ;
        RECT  6.595 -0.130 8.370 0.130 ;
        RECT  6.335 -0.130 6.595 0.400 ;
        RECT  0.385 -0.130 6.335 0.130 ;
        RECT  0.125 -0.130 0.385 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.045 2.740 10.660 3.000 ;
        RECT  8.445 2.465 9.045 3.000 ;
        RECT  4.155 2.740 8.445 3.000 ;
        RECT  3.895 2.620 4.155 3.000 ;
        RECT  0.000 2.740 3.895 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.925 1.270 10.085 2.285 ;
        RECT  8.625 2.125 9.925 2.285 ;
        RECT  9.055 1.230 9.155 1.490 ;
        RECT  8.895 0.430 9.055 1.490 ;
        RECT  8.120 0.430 8.895 0.590 ;
        RECT  8.365 0.770 8.625 2.285 ;
        RECT  8.300 1.310 8.365 1.570 ;
        RECT  7.960 0.430 8.120 2.295 ;
        RECT  7.395 0.430 7.960 0.590 ;
        RECT  7.685 2.135 7.960 2.295 ;
        RECT  7.620 0.770 7.780 1.490 ;
        RECT  7.525 2.135 7.685 2.395 ;
        RECT  7.480 1.330 7.620 1.490 ;
        RECT  7.340 1.330 7.480 1.930 ;
        RECT  7.235 0.430 7.395 0.785 ;
        RECT  7.180 1.330 7.340 2.545 ;
        RECT  6.070 0.990 7.280 1.150 ;
        RECT  6.170 1.330 7.180 1.490 ;
        RECT  4.700 2.385 7.180 2.545 ;
        RECT  6.755 1.670 6.915 2.205 ;
        RECT  5.155 2.045 6.755 2.205 ;
        RECT  5.990 1.705 6.445 1.865 ;
        RECT  6.000 0.690 6.070 1.150 ;
        RECT  5.990 0.325 6.000 1.150 ;
        RECT  5.830 0.325 5.990 1.865 ;
        RECT  3.170 0.325 5.830 0.485 ;
        RECT  5.450 0.665 5.610 1.535 ;
        RECT  5.350 0.665 5.450 0.825 ;
        RECT  5.155 1.375 5.450 1.535 ;
        RECT  3.310 1.035 5.240 1.195 ;
        RECT  4.995 1.375 5.155 2.205 ;
        RECT  3.780 1.375 4.995 1.535 ;
        RECT  4.540 2.280 4.700 2.545 ;
        RECT  4.290 0.665 4.550 0.855 ;
        RECT  3.655 2.280 4.540 2.440 ;
        RECT  2.780 0.695 4.290 0.855 ;
        RECT  3.495 2.280 3.655 2.545 ;
        RECT  2.970 2.385 3.495 2.545 ;
        RECT  3.150 1.035 3.310 2.165 ;
        RECT  2.970 1.035 3.150 1.195 ;
        RECT  2.810 1.545 2.970 2.545 ;
        RECT  2.780 1.545 2.810 1.705 ;
        RECT  2.620 0.695 2.780 1.705 ;
        RECT  0.670 0.355 2.630 0.515 ;
        RECT  2.470 1.905 2.630 2.545 ;
        RECT  0.945 2.385 2.470 2.545 ;
        RECT  0.930 0.735 1.950 0.895 ;
        RECT  0.785 2.245 0.945 2.545 ;
        RECT  0.670 0.735 0.930 1.075 ;
        RECT  0.605 1.785 0.830 1.945 ;
        RECT  0.505 0.915 0.670 1.075 ;
        RECT  0.505 1.785 0.605 2.560 ;
        RECT  0.345 0.915 0.505 2.560 ;
    END
END SDFFX2MTH

MACRO SDFFX4MTH
    CLASS CORE ;
    FOREIGN SDFFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.310 1.615 1.575 2.135 ;
        RECT  1.200 1.780 1.310 2.135 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.920 1.710 1.950 1.970 ;
        RECT  1.760 1.275 1.920 1.970 ;
        RECT  1.130 1.275 1.760 1.435 ;
        RECT  0.685 1.275 1.130 1.580 ;
        END
        AntennaGateArea 0.1053 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.805 1.290 10.970 1.580 ;
        RECT  10.545 0.405 10.805 2.390 ;
        END
        AntennaDiffArea 0.582 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.445 0.405 9.740 1.900 ;
        END
        AntennaDiffArea 0.582 ;
    END Q
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.100 1.065 2.360 1.580 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.040 1.740 4.525 1.900 ;
        RECT  3.750 1.740 4.040 2.065 ;
        END
        AntennaGateArea 0.0923 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 -0.130 11.480 0.130 ;
        RECT  11.095 -0.130 11.355 0.985 ;
        RECT  10.255 -0.130 11.095 0.130 ;
        RECT  9.995 -0.130 10.255 0.985 ;
        RECT  9.000 -0.130 9.995 0.130 ;
        RECT  8.400 -0.130 9.000 0.255 ;
        RECT  6.550 -0.130 8.400 0.130 ;
        RECT  6.290 -0.130 6.550 0.485 ;
        RECT  0.385 -0.130 6.290 0.130 ;
        RECT  0.125 -0.130 0.385 0.515 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.355 2.740 11.480 3.000 ;
        RECT  11.095 1.720 11.355 3.000 ;
        RECT  10.255 2.740 11.095 3.000 ;
        RECT  9.995 2.420 10.255 3.000 ;
        RECT  9.065 2.740 9.995 3.000 ;
        RECT  8.465 2.420 9.065 3.000 ;
        RECT  4.115 2.740 8.465 3.000 ;
        RECT  3.855 2.620 4.115 3.000 ;
        RECT  0.000 2.740 3.855 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.195 1.245 10.355 2.240 ;
        RECT  8.605 2.080 10.195 2.240 ;
        RECT  9.040 1.230 9.140 1.490 ;
        RECT  8.880 0.435 9.040 1.490 ;
        RECT  8.090 0.435 8.880 0.595 ;
        RECT  8.605 0.805 8.655 0.965 ;
        RECT  8.445 0.805 8.605 2.240 ;
        RECT  8.395 0.805 8.445 1.570 ;
        RECT  8.270 1.310 8.395 1.570 ;
        RECT  7.930 0.370 8.090 2.055 ;
        RECT  7.185 0.370 7.930 0.530 ;
        RECT  7.655 1.895 7.930 2.055 ;
        RECT  7.590 0.715 7.750 1.715 ;
        RECT  7.495 1.895 7.655 2.495 ;
        RECT  6.660 0.715 7.590 0.875 ;
        RECT  7.310 1.555 7.590 1.715 ;
        RECT  7.150 1.555 7.310 2.545 ;
        RECT  6.985 1.075 7.245 1.325 ;
        RECT  4.840 2.385 7.150 2.545 ;
        RECT  6.620 1.165 6.985 1.325 ;
        RECT  6.810 1.505 6.970 2.205 ;
        RECT  5.180 2.045 6.810 2.205 ;
        RECT  6.500 0.715 6.660 0.985 ;
        RECT  6.460 1.165 6.620 1.865 ;
        RECT  6.280 0.825 6.500 0.985 ;
        RECT  5.940 1.705 6.460 1.865 ;
        RECT  6.120 0.825 6.280 1.365 ;
        RECT  5.940 0.315 6.040 0.645 ;
        RECT  5.780 0.315 5.940 1.865 ;
        RECT  3.430 0.315 5.780 0.475 ;
        RECT  5.440 0.655 5.600 1.565 ;
        RECT  4.800 0.655 5.440 0.815 ;
        RECT  5.180 1.405 5.440 1.565 ;
        RECT  5.000 1.035 5.260 1.225 ;
        RECT  5.020 1.405 5.180 2.205 ;
        RECT  4.870 1.405 5.020 1.915 ;
        RECT  3.310 1.035 5.000 1.195 ;
        RECT  4.800 1.375 4.870 1.915 ;
        RECT  4.680 2.280 4.840 2.545 ;
        RECT  4.710 1.375 4.800 1.565 ;
        RECT  3.780 1.375 4.710 1.535 ;
        RECT  3.610 2.280 4.680 2.440 ;
        RECT  4.290 0.655 4.550 0.855 ;
        RECT  2.780 0.695 4.290 0.855 ;
        RECT  3.450 2.280 3.610 2.545 ;
        RECT  2.970 2.385 3.450 2.545 ;
        RECT  3.170 0.315 3.430 0.515 ;
        RECT  3.150 1.035 3.310 2.165 ;
        RECT  2.970 1.035 3.150 1.195 ;
        RECT  2.810 1.545 2.970 2.545 ;
        RECT  2.780 1.545 2.810 1.705 ;
        RECT  2.620 0.695 2.780 1.705 ;
        RECT  0.670 0.355 2.630 0.515 ;
        RECT  2.470 1.905 2.630 2.545 ;
        RECT  0.945 2.385 2.470 2.545 ;
        RECT  0.880 0.695 1.950 0.855 ;
        RECT  0.785 2.245 0.945 2.545 ;
        RECT  0.625 0.695 0.880 1.075 ;
        RECT  0.505 1.785 0.830 1.945 ;
        RECT  0.505 0.915 0.625 1.075 ;
        RECT  0.505 2.400 0.605 2.560 ;
        RECT  0.345 0.915 0.505 2.560 ;
    END
END SDFFX4MTH

MACRO SEDFFHQX1MTH
    CLASS CORE ;
    FOREIGN SEDFFHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.990 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.150 1.180 1.685 ;
        RECT  0.855 1.425 0.920 1.685 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.600 0.920 5.250 1.080 ;
        RECT  4.440 0.310 4.600 1.080 ;
        RECT  1.315 0.310 4.440 0.470 ;
        RECT  1.155 0.310 1.315 0.660 ;
        RECT  0.720 0.500 1.155 0.660 ;
        RECT  0.540 0.500 0.720 1.215 ;
        RECT  0.510 0.880 0.540 1.215 ;
        RECT  0.445 0.955 0.510 1.215 ;
        END
        AntennaGateArea 0.1469 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.630 0.590 15.890 2.035 ;
        RECT  15.605 0.590 15.630 0.850 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.520 1.150 5.680 1.420 ;
        RECT  5.270 1.260 5.520 1.420 ;
        RECT  4.980 1.260 5.270 1.540 ;
        RECT  4.265 1.260 4.980 1.420 ;
        RECT  4.105 1.130 4.265 1.420 ;
        END
        AntennaGateArea 0.1235 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.835 1.330 3.015 1.730 ;
        RECT  2.520 1.330 2.835 1.540 ;
        END
        AntennaGateArea 0.1131 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.925 0.920 8.960 1.170 ;
        RECT  8.585 0.680 8.925 1.170 ;
        END
        AntennaGateArea 0.1365 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.355 -0.130 15.990 0.130 ;
        RECT  15.095 -0.130 15.355 0.880 ;
        RECT  15.065 -0.130 15.095 0.300 ;
        RECT  14.740 -0.130 15.065 0.130 ;
        RECT  14.140 -0.130 14.740 0.300 ;
        RECT  12.145 -0.130 14.140 0.130 ;
        RECT  11.985 -0.130 12.145 0.300 ;
        RECT  7.565 -0.130 11.985 0.130 ;
        RECT  7.305 -0.130 7.565 0.300 ;
        RECT  5.965 -0.130 7.305 0.130 ;
        RECT  5.705 -0.130 5.965 0.300 ;
        RECT  5.040 -0.130 5.705 0.130 ;
        RECT  4.780 -0.130 5.040 0.300 ;
        RECT  0.815 -0.130 4.780 0.130 ;
        RECT  0.215 -0.130 0.815 0.300 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.545 2.740 15.990 3.000 ;
        RECT  14.605 2.570 15.545 3.000 ;
        RECT  7.745 2.740 14.605 3.000 ;
        RECT  7.145 2.620 7.745 3.000 ;
        RECT  5.625 2.740 7.145 3.000 ;
        RECT  5.025 2.280 5.625 3.000 ;
        RECT  4.155 2.740 5.025 3.000 ;
        RECT  3.895 2.620 4.155 3.000 ;
        RECT  0.845 2.740 3.895 3.000 ;
        RECT  0.245 2.570 0.845 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.235 1.130 15.285 1.390 ;
        RECT  15.075 1.130 15.235 2.215 ;
        RECT  15.025 1.130 15.075 1.390 ;
        RECT  14.490 2.055 15.075 2.215 ;
        RECT  14.685 0.615 14.845 1.815 ;
        RECT  14.575 0.615 14.685 0.875 ;
        RECT  13.960 1.180 14.685 1.340 ;
        RECT  14.330 1.715 14.490 2.215 ;
        RECT  13.615 1.715 14.330 1.875 ;
        RECT  14.075 2.400 14.175 2.560 ;
        RECT  13.915 2.060 14.075 2.560 ;
        RECT  13.800 0.310 13.960 1.340 ;
        RECT  13.275 2.060 13.915 2.220 ;
        RECT  12.485 0.310 13.800 0.470 ;
        RECT  10.785 2.400 13.635 2.560 ;
        RECT  13.455 0.650 13.615 1.875 ;
        RECT  13.175 0.650 13.455 0.810 ;
        RECT  13.115 0.990 13.275 2.220 ;
        RECT  11.125 2.060 13.115 2.220 ;
        RECT  12.775 0.650 12.935 1.850 ;
        RECT  12.665 0.650 12.775 0.980 ;
        RECT  12.115 0.820 12.665 0.980 ;
        RECT  12.485 1.180 12.595 1.440 ;
        RECT  12.325 0.310 12.485 0.640 ;
        RECT  12.325 1.180 12.485 1.780 ;
        RECT  11.805 0.480 12.325 0.640 ;
        RECT  11.775 1.620 12.325 1.780 ;
        RECT  11.955 0.820 12.115 1.265 ;
        RECT  11.645 0.310 11.805 0.640 ;
        RECT  11.615 0.820 11.775 1.780 ;
        RECT  7.910 0.310 11.645 0.470 ;
        RECT  11.465 0.820 11.615 0.980 ;
        RECT  11.465 1.620 11.615 1.780 ;
        RECT  11.205 0.650 11.465 0.980 ;
        RECT  11.305 1.620 11.465 1.880 ;
        RECT  11.125 1.160 11.435 1.420 ;
        RECT  11.025 1.160 11.125 2.220 ;
        RECT  10.965 0.650 11.025 2.220 ;
        RECT  10.865 0.650 10.965 1.320 ;
        RECT  10.035 0.650 10.865 0.810 ;
        RECT  10.685 2.055 10.785 2.560 ;
        RECT  10.625 0.990 10.685 2.560 ;
        RECT  10.525 0.990 10.625 2.220 ;
        RECT  10.425 0.990 10.525 1.150 ;
        RECT  8.420 2.060 10.525 2.220 ;
        RECT  8.085 2.400 10.400 2.560 ;
        RECT  10.035 1.335 10.205 1.495 ;
        RECT  9.875 0.650 10.035 1.875 ;
        RECT  9.675 0.650 9.875 0.810 ;
        RECT  8.860 1.715 9.875 1.875 ;
        RECT  9.410 1.250 9.610 1.510 ;
        RECT  9.250 0.650 9.410 1.510 ;
        RECT  9.150 0.650 9.250 0.810 ;
        RECT  8.360 1.350 9.250 1.510 ;
        RECT  8.600 1.690 8.860 1.875 ;
        RECT  8.260 1.925 8.420 2.220 ;
        RECT  8.250 0.655 8.405 0.815 ;
        RECT  8.200 1.350 8.360 1.745 ;
        RECT  7.920 1.925 8.260 2.085 ;
        RECT  8.090 0.655 8.250 1.170 ;
        RECT  8.100 1.585 8.200 1.745 ;
        RECT  7.920 1.010 8.090 1.170 ;
        RECT  7.925 2.270 8.085 2.560 ;
        RECT  6.900 2.270 7.925 2.430 ;
        RECT  7.760 1.010 7.920 2.085 ;
        RECT  7.750 0.310 7.910 0.825 ;
        RECT  7.580 0.665 7.750 0.825 ;
        RECT  7.420 0.665 7.580 1.440 ;
        RECT  6.935 0.485 7.095 1.830 ;
        RECT  6.785 0.485 6.935 0.745 ;
        RECT  6.900 1.570 6.935 1.830 ;
        RECT  6.740 1.570 6.900 2.560 ;
        RECT  6.560 1.230 6.755 1.390 ;
        RECT  5.965 2.400 6.740 2.560 ;
        RECT  6.400 0.500 6.560 2.220 ;
        RECT  6.325 0.500 6.400 0.760 ;
        RECT  6.210 2.060 6.400 2.220 ;
        RECT  6.065 0.965 6.220 1.565 ;
        RECT  5.905 0.550 6.065 1.760 ;
        RECT  5.805 1.940 5.965 2.560 ;
        RECT  5.245 0.550 5.905 0.710 ;
        RECT  5.640 1.600 5.905 1.760 ;
        RECT  3.225 1.940 5.805 2.100 ;
        RECT  3.675 2.280 4.785 2.440 ;
        RECT  3.925 1.600 4.575 1.760 ;
        RECT  3.925 0.650 4.115 0.810 ;
        RECT  3.765 0.650 3.925 1.760 ;
        RECT  3.535 1.095 3.765 1.355 ;
        RECT  3.515 2.280 3.675 2.560 ;
        RECT  3.355 1.570 3.585 1.730 ;
        RECT  3.355 0.650 3.575 0.910 ;
        RECT  1.305 2.400 3.515 2.560 ;
        RECT  3.195 0.650 3.355 1.730 ;
        RECT  3.065 1.940 3.225 2.220 ;
        RECT  2.335 0.990 3.195 1.150 ;
        RECT  1.695 2.060 3.065 2.220 ;
        RECT  2.260 1.720 2.655 1.880 ;
        RECT  1.995 0.650 2.440 0.810 ;
        RECT  2.175 0.990 2.335 1.250 ;
        RECT  2.100 1.430 2.260 1.880 ;
        RECT  1.995 1.430 2.100 1.590 ;
        RECT  1.835 0.650 1.995 1.590 ;
        RECT  1.655 1.725 1.695 2.220 ;
        RECT  1.495 0.675 1.655 2.220 ;
        RECT  1.145 1.895 1.305 2.560 ;
        RECT  0.385 1.895 1.145 2.055 ;
        RECT  0.265 1.795 0.385 2.055 ;
        RECT  0.265 0.550 0.335 0.810 ;
        RECT  0.105 0.550 0.265 2.055 ;
    END
END SEDFFHQX1MTH

MACRO SEDFFHQX2MTH
    CLASS CORE ;
    FOREIGN SEDFFHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.990 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.150 1.180 1.700 ;
        RECT  0.855 1.440 0.920 1.700 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.595 0.920 5.250 1.080 ;
        RECT  4.435 0.310 4.595 1.080 ;
        RECT  1.305 0.310 4.435 0.470 ;
        RECT  1.145 0.310 1.305 0.660 ;
        RECT  0.740 0.500 1.145 0.660 ;
        RECT  0.550 0.500 0.740 1.230 ;
        RECT  0.510 0.880 0.550 1.230 ;
        RECT  0.445 0.970 0.510 1.230 ;
        END
        AntennaGateArea 0.1469 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  15.630 0.390 15.890 2.425 ;
        RECT  15.605 0.390 15.630 0.990 ;
        RECT  15.605 1.825 15.630 2.425 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.520 1.150 5.680 1.420 ;
        RECT  5.270 1.260 5.520 1.420 ;
        RECT  4.980 1.260 5.270 1.540 ;
        RECT  4.255 1.260 4.980 1.420 ;
        RECT  4.095 1.130 4.255 1.420 ;
        END
        AntennaGateArea 0.117 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.825 1.330 3.015 1.730 ;
        RECT  2.520 1.330 2.825 1.540 ;
        END
        AntennaGateArea 0.0923 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.925 0.920 8.960 1.170 ;
        RECT  8.530 0.680 8.925 1.170 ;
        END
        AntennaGateArea 0.1443 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.355 -0.130 15.990 0.130 ;
        RECT  15.095 -0.130 15.355 0.945 ;
        RECT  14.915 -0.130 15.095 0.130 ;
        RECT  14.315 -0.130 14.915 0.300 ;
        RECT  12.105 -0.130 14.315 0.130 ;
        RECT  11.945 -0.130 12.105 0.300 ;
        RECT  7.565 -0.130 11.945 0.130 ;
        RECT  7.305 -0.130 7.565 0.300 ;
        RECT  5.965 -0.130 7.305 0.130 ;
        RECT  5.705 -0.130 5.965 0.300 ;
        RECT  5.035 -0.130 5.705 0.130 ;
        RECT  4.775 -0.130 5.035 0.300 ;
        RECT  0.965 -0.130 4.775 0.130 ;
        RECT  0.365 -0.130 0.965 0.300 ;
        RECT  0.000 -0.130 0.365 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.325 2.740 15.990 3.000 ;
        RECT  14.385 2.570 15.325 3.000 ;
        RECT  7.755 2.740 14.385 3.000 ;
        RECT  7.155 2.620 7.755 3.000 ;
        RECT  5.625 2.740 7.155 3.000 ;
        RECT  5.025 2.280 5.625 3.000 ;
        RECT  4.360 2.740 5.025 3.000 ;
        RECT  3.760 2.620 4.360 3.000 ;
        RECT  0.845 2.740 3.760 3.000 ;
        RECT  0.245 2.570 0.845 3.000 ;
        RECT  0.000 2.740 0.245 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.085 1.205 15.445 1.465 ;
        RECT  14.925 1.205 15.085 2.220 ;
        RECT  14.365 2.060 14.925 2.220 ;
        RECT  14.715 0.695 14.775 0.955 ;
        RECT  14.555 0.695 14.715 1.875 ;
        RECT  14.025 1.080 14.555 1.240 ;
        RECT  14.205 1.420 14.365 2.220 ;
        RECT  13.685 1.420 14.205 1.580 ;
        RECT  13.865 0.310 14.025 1.240 ;
        RECT  13.865 1.760 14.025 2.220 ;
        RECT  12.445 0.310 13.865 0.470 ;
        RECT  13.245 2.060 13.865 2.220 ;
        RECT  10.885 2.400 13.690 2.560 ;
        RECT  13.525 0.650 13.685 1.875 ;
        RECT  13.135 0.650 13.525 0.810 ;
        RECT  13.425 1.715 13.525 1.875 ;
        RECT  13.245 1.035 13.345 1.195 ;
        RECT  13.085 1.035 13.245 2.220 ;
        RECT  11.225 2.060 13.085 2.220 ;
        RECT  12.745 0.650 12.905 1.880 ;
        RECT  12.625 0.650 12.745 0.980 ;
        RECT  12.645 1.720 12.745 1.880 ;
        RECT  12.085 0.820 12.625 0.980 ;
        RECT  12.465 1.195 12.565 1.455 ;
        RECT  12.305 1.195 12.465 1.780 ;
        RECT  12.285 0.310 12.445 0.640 ;
        RECT  11.745 1.620 12.305 1.780 ;
        RECT  11.765 0.480 12.285 0.640 ;
        RECT  11.925 0.820 12.085 1.305 ;
        RECT  11.605 0.310 11.765 0.640 ;
        RECT  11.585 0.820 11.745 1.780 ;
        RECT  7.910 0.310 11.605 0.470 ;
        RECT  11.425 0.820 11.585 0.980 ;
        RECT  11.565 1.620 11.585 1.780 ;
        RECT  11.405 1.620 11.565 1.880 ;
        RECT  11.165 0.650 11.425 0.980 ;
        RECT  11.225 1.160 11.405 1.420 ;
        RECT  11.065 1.160 11.225 2.220 ;
        RECT  10.980 1.160 11.065 1.420 ;
        RECT  10.820 0.650 10.980 1.420 ;
        RECT  10.725 2.060 10.885 2.560 ;
        RECT  10.015 0.650 10.820 0.810 ;
        RECT  10.640 2.060 10.725 2.220 ;
        RECT  10.480 1.020 10.640 2.220 ;
        RECT  8.085 2.400 10.545 2.560 ;
        RECT  10.380 1.020 10.480 1.180 ;
        RECT  8.425 2.060 10.480 2.220 ;
        RECT  9.855 0.650 10.015 1.875 ;
        RECT  9.615 0.650 9.855 0.810 ;
        RECT  8.865 1.715 9.855 1.875 ;
        RECT  9.365 1.180 9.585 1.440 ;
        RECT  9.205 0.650 9.365 1.510 ;
        RECT  9.105 0.650 9.205 0.810 ;
        RECT  8.335 1.350 9.205 1.510 ;
        RECT  8.605 1.690 8.865 1.875 ;
        RECT  8.265 1.925 8.425 2.220 ;
        RECT  8.250 0.650 8.350 0.810 ;
        RECT  8.175 1.350 8.335 1.745 ;
        RECT  7.895 1.925 8.265 2.085 ;
        RECT  8.090 0.650 8.250 1.070 ;
        RECT  8.075 1.585 8.175 1.745 ;
        RECT  7.895 0.910 8.090 1.070 ;
        RECT  7.925 2.270 8.085 2.560 ;
        RECT  6.825 2.270 7.925 2.430 ;
        RECT  7.750 0.310 7.910 0.720 ;
        RECT  7.735 0.910 7.895 2.085 ;
        RECT  7.555 0.560 7.750 0.720 ;
        RECT  7.395 0.560 7.555 1.440 ;
        RECT  6.935 0.485 7.095 1.775 ;
        RECT  6.835 0.485 6.935 0.745 ;
        RECT  6.825 1.615 6.935 1.775 ;
        RECT  6.665 1.615 6.825 2.560 ;
        RECT  6.610 1.190 6.755 1.435 ;
        RECT  5.965 2.400 6.665 2.560 ;
        RECT  6.485 0.550 6.610 1.435 ;
        RECT  6.450 0.550 6.485 2.220 ;
        RECT  6.275 0.550 6.450 0.710 ;
        RECT  6.325 1.275 6.450 2.220 ;
        RECT  6.210 2.060 6.325 2.220 ;
        RECT  6.065 0.920 6.270 1.080 ;
        RECT  5.905 0.550 6.065 1.760 ;
        RECT  5.805 1.940 5.965 2.560 ;
        RECT  5.245 0.550 5.905 0.710 ;
        RECT  5.640 1.600 5.905 1.760 ;
        RECT  3.185 1.940 5.805 2.100 ;
        RECT  3.555 2.280 4.785 2.440 ;
        RECT  3.915 1.600 4.575 1.760 ;
        RECT  3.915 0.650 4.105 0.810 ;
        RECT  3.755 0.650 3.915 1.760 ;
        RECT  3.565 1.040 3.755 1.300 ;
        RECT  3.385 0.650 3.575 0.810 ;
        RECT  3.385 1.570 3.575 1.730 ;
        RECT  3.395 2.280 3.555 2.560 ;
        RECT  1.260 2.400 3.395 2.560 ;
        RECT  3.225 0.650 3.385 1.730 ;
        RECT  2.335 0.990 3.225 1.150 ;
        RECT  3.025 1.940 3.185 2.220 ;
        RECT  1.745 2.060 3.025 2.220 ;
        RECT  2.260 1.720 2.645 1.880 ;
        RECT  1.995 0.650 2.525 0.810 ;
        RECT  2.175 0.990 2.335 1.250 ;
        RECT  2.100 1.430 2.260 1.880 ;
        RECT  1.995 1.430 2.100 1.590 ;
        RECT  1.835 0.650 1.995 1.590 ;
        RECT  1.655 1.775 1.745 2.220 ;
        RECT  1.485 0.675 1.655 2.220 ;
        RECT  1.100 1.910 1.260 2.560 ;
        RECT  0.385 1.910 1.100 2.070 ;
        RECT  0.265 1.810 0.385 2.070 ;
        RECT  0.265 0.555 0.335 0.815 ;
        RECT  0.105 0.555 0.265 2.070 ;
    END
END SEDFFHQX2MTH

MACRO SEDFFHQX4MTH
    CLASS CORE ;
    FOREIGN SEDFFHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.810 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.150 1.180 1.685 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.005 0.920 5.660 1.080 ;
        RECT  4.845 0.310 5.005 1.080 ;
        RECT  3.545 0.310 4.845 0.470 ;
        RECT  3.385 0.310 3.545 0.640 ;
        RECT  2.865 0.480 3.385 0.640 ;
        RECT  2.705 0.310 2.865 0.640 ;
        RECT  1.160 0.310 2.705 0.470 ;
        RECT  1.000 0.310 1.160 0.660 ;
        RECT  0.720 0.500 1.000 0.660 ;
        RECT  0.540 0.500 0.720 1.415 ;
        RECT  0.510 0.880 0.540 1.415 ;
        RECT  0.470 1.155 0.510 1.415 ;
        END
        AntennaGateArea 0.1469 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.175 1.290 16.300 1.580 ;
        RECT  15.915 0.390 16.175 2.425 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.930 1.150 6.090 1.420 ;
        RECT  5.680 1.260 5.930 1.420 ;
        RECT  5.390 1.260 5.680 1.540 ;
        RECT  4.665 1.260 5.390 1.420 ;
        RECT  4.505 1.130 4.665 1.420 ;
        END
        AntennaGateArea 0.117 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.330 3.150 1.540 ;
        END
        AntennaGateArea 0.1638 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.335 0.920 9.370 1.170 ;
        RECT  8.955 0.680 9.335 1.170 ;
        RECT  8.870 1.010 8.955 1.170 ;
        END
        AntennaGateArea 0.1859 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.685 -0.130 16.810 0.130 ;
        RECT  16.425 -0.130 16.685 0.990 ;
        RECT  15.635 -0.130 16.425 0.130 ;
        RECT  15.035 -0.130 15.635 0.300 ;
        RECT  12.565 -0.130 15.035 0.130 ;
        RECT  12.405 -0.130 12.565 0.300 ;
        RECT  7.975 -0.130 12.405 0.130 ;
        RECT  7.715 -0.130 7.975 0.300 ;
        RECT  6.375 -0.130 7.715 0.130 ;
        RECT  6.115 -0.130 6.375 0.300 ;
        RECT  5.445 -0.130 6.115 0.130 ;
        RECT  5.185 -0.130 5.445 0.300 ;
        RECT  3.205 -0.130 5.185 0.130 ;
        RECT  3.045 -0.130 3.205 0.300 ;
        RECT  0.815 -0.130 3.045 0.130 ;
        RECT  0.215 -0.130 0.815 0.300 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.685 2.740 16.810 3.000 ;
        RECT  16.425 1.825 16.685 3.000 ;
        RECT  15.635 2.740 16.425 3.000 ;
        RECT  15.035 2.570 15.635 3.000 ;
        RECT  8.155 2.740 15.035 3.000 ;
        RECT  7.555 2.620 8.155 3.000 ;
        RECT  6.035 2.740 7.555 3.000 ;
        RECT  5.435 2.280 6.035 3.000 ;
        RECT  4.770 2.740 5.435 3.000 ;
        RECT  4.510 2.620 4.770 3.000 ;
        RECT  0.965 2.740 4.510 3.000 ;
        RECT  0.365 2.570 0.965 3.000 ;
        RECT  0.000 2.740 0.365 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.425 1.205 15.585 2.365 ;
        RECT  14.815 2.205 15.425 2.365 ;
        RECT  14.995 0.765 15.155 1.945 ;
        RECT  14.785 0.765 14.995 0.925 ;
        RECT  14.655 1.420 14.815 2.365 ;
        RECT  14.625 0.310 14.785 1.195 ;
        RECT  14.405 1.420 14.655 1.580 ;
        RECT  12.905 0.310 14.625 0.470 ;
        RECT  14.305 1.760 14.465 2.220 ;
        RECT  14.245 0.650 14.405 1.580 ;
        RECT  13.655 2.060 14.305 2.220 ;
        RECT  13.525 0.650 14.245 0.810 ;
        RECT  14.095 1.420 14.245 1.580 ;
        RECT  13.935 1.420 14.095 1.875 ;
        RECT  11.295 2.400 14.085 2.560 ;
        RECT  13.655 1.020 14.045 1.180 ;
        RECT  13.835 1.715 13.935 1.875 ;
        RECT  13.495 1.020 13.655 2.220 ;
        RECT  11.635 2.060 13.495 2.220 ;
        RECT  13.155 0.745 13.315 1.880 ;
        RECT  13.065 0.745 13.155 1.005 ;
        RECT  13.055 1.720 13.155 1.880 ;
        RECT  12.495 0.820 13.065 0.980 ;
        RECT  12.875 1.195 12.975 1.455 ;
        RECT  12.745 0.310 12.905 0.640 ;
        RECT  12.715 1.195 12.875 1.780 ;
        RECT  12.175 0.480 12.745 0.640 ;
        RECT  12.155 1.620 12.715 1.780 ;
        RECT  12.335 0.820 12.495 1.375 ;
        RECT  12.015 0.310 12.175 0.640 ;
        RECT  11.995 0.820 12.155 1.780 ;
        RECT  8.320 0.310 12.015 0.470 ;
        RECT  11.835 0.820 11.995 0.980 ;
        RECT  11.975 1.620 11.995 1.780 ;
        RECT  11.815 1.620 11.975 1.880 ;
        RECT  11.575 0.650 11.835 0.980 ;
        RECT  11.635 1.160 11.815 1.420 ;
        RECT  11.475 1.160 11.635 2.220 ;
        RECT  11.390 1.160 11.475 1.420 ;
        RECT  11.230 0.650 11.390 1.420 ;
        RECT  11.135 2.060 11.295 2.560 ;
        RECT  10.425 0.650 11.230 0.810 ;
        RECT  10.950 2.060 11.135 2.220 ;
        RECT  10.950 0.990 11.050 1.150 ;
        RECT  8.495 2.400 10.955 2.560 ;
        RECT  10.790 0.990 10.950 2.220 ;
        RECT  8.835 2.060 10.790 2.220 ;
        RECT  10.265 0.650 10.425 1.875 ;
        RECT  10.025 0.650 10.265 0.810 ;
        RECT  9.275 1.715 10.265 1.875 ;
        RECT  9.775 1.180 9.995 1.440 ;
        RECT  9.615 0.650 9.775 1.510 ;
        RECT  9.515 0.650 9.615 0.810 ;
        RECT  8.745 1.350 9.615 1.510 ;
        RECT  9.015 1.690 9.275 1.875 ;
        RECT  8.675 1.925 8.835 2.220 ;
        RECT  8.675 0.650 8.775 0.810 ;
        RECT  8.585 1.350 8.745 1.730 ;
        RECT  8.515 0.650 8.675 1.070 ;
        RECT  8.305 1.925 8.675 2.085 ;
        RECT  8.485 1.570 8.585 1.730 ;
        RECT  8.305 0.910 8.515 1.070 ;
        RECT  8.335 2.270 8.495 2.560 ;
        RECT  7.235 2.270 8.335 2.430 ;
        RECT  8.160 0.310 8.320 0.720 ;
        RECT  8.145 0.910 8.305 2.085 ;
        RECT  7.965 0.560 8.160 0.720 ;
        RECT  7.805 0.560 7.965 1.460 ;
        RECT  7.700 1.200 7.805 1.460 ;
        RECT  7.345 0.520 7.505 2.090 ;
        RECT  7.245 0.520 7.345 0.780 ;
        RECT  7.235 1.930 7.345 2.090 ;
        RECT  7.075 1.930 7.235 2.560 ;
        RECT  7.020 1.515 7.165 1.750 ;
        RECT  6.375 2.400 7.075 2.560 ;
        RECT  6.895 0.550 7.020 1.750 ;
        RECT  6.860 0.550 6.895 2.220 ;
        RECT  6.685 0.550 6.860 0.710 ;
        RECT  6.735 1.560 6.860 2.220 ;
        RECT  6.620 2.060 6.735 2.220 ;
        RECT  6.475 0.940 6.680 1.100 ;
        RECT  6.315 0.550 6.475 1.760 ;
        RECT  6.215 1.940 6.375 2.560 ;
        RECT  5.655 0.550 6.315 0.710 ;
        RECT  6.050 1.600 6.315 1.760 ;
        RECT  3.575 1.940 6.215 2.100 ;
        RECT  4.295 2.280 5.195 2.440 ;
        RECT  4.325 1.600 4.985 1.760 ;
        RECT  4.325 0.650 4.515 0.810 ;
        RECT  4.165 0.650 4.325 1.760 ;
        RECT  4.135 2.280 4.295 2.560 ;
        RECT  4.025 1.130 4.165 1.390 ;
        RECT  1.315 2.400 4.135 2.560 ;
        RECT  3.845 0.650 3.985 0.950 ;
        RECT  3.845 1.570 3.945 1.730 ;
        RECT  3.725 0.650 3.845 1.730 ;
        RECT  3.685 0.760 3.725 1.730 ;
        RECT  2.335 0.990 3.685 1.150 ;
        RECT  3.415 1.940 3.575 2.220 ;
        RECT  1.865 2.060 3.415 2.220 ;
        RECT  2.305 1.720 3.035 1.880 ;
        RECT  1.995 0.650 2.525 0.810 ;
        RECT  2.175 0.990 2.335 1.255 ;
        RECT  2.145 1.435 2.305 1.880 ;
        RECT  1.995 1.435 2.145 1.595 ;
        RECT  1.835 0.650 1.995 1.595 ;
        RECT  1.655 1.775 1.865 2.220 ;
        RECT  1.495 0.675 1.655 2.220 ;
        RECT  1.155 1.895 1.315 2.560 ;
        RECT  0.385 1.895 1.155 2.055 ;
        RECT  0.270 1.795 0.385 2.055 ;
        RECT  0.270 0.555 0.335 0.815 ;
        RECT  0.110 0.555 0.270 2.055 ;
    END
END SEDFFHQX4MTH

MACRO SEDFFHQX8MTH
    CLASS CORE ;
    FOREIGN SEDFFHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.040 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.915 1.150 1.180 1.685 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.005 0.920 5.660 1.080 ;
        RECT  4.845 0.310 5.005 1.080 ;
        RECT  3.545 0.310 4.845 0.470 ;
        RECT  3.385 0.310 3.545 0.640 ;
        RECT  2.865 0.480 3.385 0.640 ;
        RECT  2.705 0.310 2.865 0.640 ;
        RECT  1.160 0.310 2.705 0.470 ;
        RECT  1.000 0.310 1.160 0.660 ;
        RECT  0.720 0.500 1.000 0.660 ;
        RECT  0.540 0.500 0.720 1.415 ;
        RECT  0.510 0.880 0.540 1.415 ;
        RECT  0.470 1.155 0.510 1.415 ;
        END
        AntennaGateArea 0.1469 ;
    END SE
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.145 0.390 17.405 2.425 ;
        RECT  16.385 1.290 17.145 1.580 ;
        RECT  16.125 0.390 16.385 2.425 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.930 1.150 6.090 1.420 ;
        RECT  5.680 1.260 5.930 1.420 ;
        RECT  5.390 1.260 5.680 1.540 ;
        RECT  4.665 1.260 5.390 1.420 ;
        RECT  4.505 1.130 4.665 1.420 ;
        END
        AntennaGateArea 0.117 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.330 3.150 1.540 ;
        END
        AntennaGateArea 0.1638 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.335 0.920 9.370 1.170 ;
        RECT  8.955 0.680 9.335 1.170 ;
        RECT  8.870 1.010 8.955 1.170 ;
        END
        AntennaGateArea 0.1859 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.915 -0.130 18.040 0.130 ;
        RECT  17.655 -0.130 17.915 0.990 ;
        RECT  16.895 -0.130 17.655 0.130 ;
        RECT  16.635 -0.130 16.895 0.990 ;
        RECT  15.840 -0.130 16.635 0.130 ;
        RECT  15.560 -0.130 15.840 0.990 ;
        RECT  14.965 -0.130 15.560 0.300 ;
        RECT  12.565 -0.130 14.965 0.130 ;
        RECT  12.405 -0.130 12.565 0.300 ;
        RECT  7.975 -0.130 12.405 0.130 ;
        RECT  7.715 -0.130 7.975 0.300 ;
        RECT  6.375 -0.130 7.715 0.130 ;
        RECT  6.115 -0.130 6.375 0.300 ;
        RECT  5.445 -0.130 6.115 0.130 ;
        RECT  5.185 -0.130 5.445 0.300 ;
        RECT  3.205 -0.130 5.185 0.130 ;
        RECT  3.045 -0.130 3.205 0.300 ;
        RECT  0.815 -0.130 3.045 0.130 ;
        RECT  0.215 -0.130 0.815 0.300 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.915 2.740 18.040 3.000 ;
        RECT  17.655 1.825 17.915 3.000 ;
        RECT  16.895 2.740 17.655 3.000 ;
        RECT  16.635 1.825 16.895 3.000 ;
        RECT  15.635 2.740 16.635 3.000 ;
        RECT  15.035 2.570 15.635 3.000 ;
        RECT  8.155 2.740 15.035 3.000 ;
        RECT  7.555 2.620 8.155 3.000 ;
        RECT  6.035 2.740 7.555 3.000 ;
        RECT  5.435 2.280 6.035 3.000 ;
        RECT  4.770 2.740 5.435 3.000 ;
        RECT  4.510 2.620 4.770 3.000 ;
        RECT  0.965 2.740 4.510 3.000 ;
        RECT  0.365 2.570 0.965 3.000 ;
        RECT  0.000 2.740 0.365 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.620 1.205 15.945 1.465 ;
        RECT  15.460 1.205 15.620 2.365 ;
        RECT  15.345 1.205 15.460 1.465 ;
        RECT  14.815 2.205 15.460 2.365 ;
        RECT  14.995 0.765 15.155 1.945 ;
        RECT  14.785 0.765 14.995 1.195 ;
        RECT  14.655 1.420 14.815 2.365 ;
        RECT  14.625 0.310 14.785 1.195 ;
        RECT  14.405 1.420 14.655 1.580 ;
        RECT  12.905 0.310 14.625 0.470 ;
        RECT  14.305 1.760 14.465 2.220 ;
        RECT  14.245 0.650 14.405 1.580 ;
        RECT  13.655 2.060 14.305 2.220 ;
        RECT  13.525 0.650 14.245 0.810 ;
        RECT  14.095 1.420 14.245 1.580 ;
        RECT  13.935 1.420 14.095 1.875 ;
        RECT  11.295 2.400 14.085 2.560 ;
        RECT  13.655 1.020 14.045 1.180 ;
        RECT  13.835 1.715 13.935 1.875 ;
        RECT  13.495 1.020 13.655 2.220 ;
        RECT  11.635 2.060 13.495 2.220 ;
        RECT  13.155 0.745 13.315 1.880 ;
        RECT  13.065 0.745 13.155 1.005 ;
        RECT  13.055 1.720 13.155 1.880 ;
        RECT  12.495 0.820 13.065 0.980 ;
        RECT  12.875 1.195 12.975 1.455 ;
        RECT  12.745 0.310 12.905 0.640 ;
        RECT  12.715 1.195 12.875 1.780 ;
        RECT  12.175 0.480 12.745 0.640 ;
        RECT  12.155 1.620 12.715 1.780 ;
        RECT  12.335 0.820 12.495 1.375 ;
        RECT  12.015 0.310 12.175 0.640 ;
        RECT  11.995 0.820 12.155 1.780 ;
        RECT  8.320 0.310 12.015 0.470 ;
        RECT  11.835 0.820 11.995 0.980 ;
        RECT  11.975 1.620 11.995 1.780 ;
        RECT  11.815 1.620 11.975 1.880 ;
        RECT  11.575 0.650 11.835 0.980 ;
        RECT  11.635 1.160 11.815 1.420 ;
        RECT  11.475 1.160 11.635 2.220 ;
        RECT  11.390 1.160 11.475 1.420 ;
        RECT  11.230 0.650 11.390 1.420 ;
        RECT  11.135 2.060 11.295 2.560 ;
        RECT  10.425 0.650 11.230 0.810 ;
        RECT  10.950 2.060 11.135 2.220 ;
        RECT  10.950 0.990 11.050 1.150 ;
        RECT  8.495 2.400 10.955 2.560 ;
        RECT  10.790 0.990 10.950 2.220 ;
        RECT  8.835 2.060 10.790 2.220 ;
        RECT  10.265 0.650 10.425 1.875 ;
        RECT  10.025 0.650 10.265 0.810 ;
        RECT  9.275 1.715 10.265 1.875 ;
        RECT  9.775 1.180 9.995 1.440 ;
        RECT  9.615 0.650 9.775 1.510 ;
        RECT  9.515 0.650 9.615 0.810 ;
        RECT  8.745 1.350 9.615 1.510 ;
        RECT  9.015 1.690 9.275 1.875 ;
        RECT  8.675 1.925 8.835 2.220 ;
        RECT  8.675 0.650 8.775 0.810 ;
        RECT  8.585 1.350 8.745 1.730 ;
        RECT  8.515 0.650 8.675 1.070 ;
        RECT  8.305 1.925 8.675 2.085 ;
        RECT  8.485 1.570 8.585 1.730 ;
        RECT  8.305 0.910 8.515 1.070 ;
        RECT  8.335 2.270 8.495 2.560 ;
        RECT  7.235 2.270 8.335 2.430 ;
        RECT  8.160 0.310 8.320 0.720 ;
        RECT  8.145 0.910 8.305 2.085 ;
        RECT  7.965 0.560 8.160 0.720 ;
        RECT  7.805 0.560 7.965 1.460 ;
        RECT  7.700 1.200 7.805 1.460 ;
        RECT  7.345 0.520 7.505 2.090 ;
        RECT  7.245 0.520 7.345 0.780 ;
        RECT  7.235 1.930 7.345 2.090 ;
        RECT  7.075 1.930 7.235 2.560 ;
        RECT  7.020 1.515 7.165 1.750 ;
        RECT  6.375 2.400 7.075 2.560 ;
        RECT  6.895 0.550 7.020 1.750 ;
        RECT  6.860 0.550 6.895 2.220 ;
        RECT  6.685 0.550 6.860 0.710 ;
        RECT  6.735 1.560 6.860 2.220 ;
        RECT  6.620 2.060 6.735 2.220 ;
        RECT  6.475 0.940 6.680 1.100 ;
        RECT  6.315 0.550 6.475 1.760 ;
        RECT  6.215 1.940 6.375 2.560 ;
        RECT  5.655 0.550 6.315 0.710 ;
        RECT  6.050 1.600 6.315 1.760 ;
        RECT  3.575 1.940 6.215 2.100 ;
        RECT  4.295 2.280 5.195 2.440 ;
        RECT  4.325 1.600 4.985 1.760 ;
        RECT  4.325 0.650 4.515 0.810 ;
        RECT  4.165 0.650 4.325 1.760 ;
        RECT  4.135 2.280 4.295 2.560 ;
        RECT  4.025 1.130 4.165 1.390 ;
        RECT  1.315 2.400 4.135 2.560 ;
        RECT  3.845 0.650 3.985 0.950 ;
        RECT  3.845 1.570 3.945 1.730 ;
        RECT  3.725 0.650 3.845 1.730 ;
        RECT  3.685 0.760 3.725 1.730 ;
        RECT  2.335 0.990 3.685 1.150 ;
        RECT  3.415 1.940 3.575 2.220 ;
        RECT  1.865 2.060 3.415 2.220 ;
        RECT  2.305 1.720 3.035 1.880 ;
        RECT  1.995 0.650 2.525 0.810 ;
        RECT  2.175 0.990 2.335 1.250 ;
        RECT  2.145 1.430 2.305 1.880 ;
        RECT  1.995 1.430 2.145 1.590 ;
        RECT  1.835 0.650 1.995 1.590 ;
        RECT  1.655 1.775 1.865 2.220 ;
        RECT  1.495 0.675 1.655 2.220 ;
        RECT  1.155 1.895 1.315 2.560 ;
        RECT  0.385 1.895 1.155 2.055 ;
        RECT  0.270 1.795 0.385 2.055 ;
        RECT  0.270 0.555 0.335 0.815 ;
        RECT  0.110 0.555 0.270 2.055 ;
    END
END SEDFFHQX8MTH

MACRO SEDFFTRX1MTH
    CLASS CORE ;
    FOREIGN SEDFFTRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.860 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.200 2.075 1.460 ;
        RECT  1.740 1.200 1.975 1.720 ;
        END
        AntennaGateArea 0.052 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 1.175 1.540 1.720 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.790 0.440 1.170 ;
        END
        AntennaGateArea 0.0624 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.730 0.815 17.940 2.080 ;
        RECT  17.535 0.815 17.730 0.975 ;
        RECT  17.555 1.820 17.730 2.080 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.605 0.720 18.765 2.060 ;
        RECT  18.475 0.720 18.605 0.980 ;
        RECT  18.495 1.670 18.605 2.060 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.260 1.330 7.730 1.575 ;
        RECT  7.160 1.330 7.260 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 1.190 4.980 1.450 ;
        RECT  4.520 1.190 4.910 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 1.205 9.185 1.725 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.365 -0.130 18.860 0.130 ;
        RECT  17.425 -0.130 18.365 0.250 ;
        RECT  14.765 -0.130 17.425 0.130 ;
        RECT  14.605 -0.130 14.765 0.915 ;
        RECT  12.835 -0.130 14.605 0.130 ;
        RECT  12.675 -0.130 12.835 0.645 ;
        RECT  11.135 -0.130 12.675 0.130 ;
        RECT  10.915 -0.130 11.135 1.025 ;
        RECT  9.895 -0.130 10.915 0.130 ;
        RECT  8.955 -0.130 9.895 0.250 ;
        RECT  5.110 -0.130 8.955 0.130 ;
        RECT  4.510 -0.130 5.110 0.250 ;
        RECT  1.450 -0.130 4.510 0.130 ;
        RECT  1.190 -0.130 1.450 0.305 ;
        RECT  0.725 -0.130 1.190 0.130 ;
        RECT  0.125 -0.130 0.725 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.185 2.740 18.860 3.000 ;
        RECT  17.585 2.620 18.185 3.000 ;
        RECT  17.225 2.740 17.585 3.000 ;
        RECT  16.625 2.620 17.225 3.000 ;
        RECT  12.935 2.740 16.625 3.000 ;
        RECT  12.675 2.620 12.935 3.000 ;
        RECT  10.305 2.740 12.675 3.000 ;
        RECT  10.045 2.295 10.305 3.000 ;
        RECT  8.845 2.740 10.045 3.000 ;
        RECT  8.685 2.245 8.845 3.000 ;
        RECT  1.245 2.740 8.685 3.000 ;
        RECT  0.985 2.620 1.245 3.000 ;
        RECT  0.000 2.740 0.985 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.280 1.205 18.405 1.465 ;
        RECT  18.120 0.475 18.280 2.440 ;
        RECT  17.235 0.475 18.120 0.635 ;
        RECT  17.235 2.280 18.120 2.440 ;
        RECT  16.895 1.205 17.455 1.465 ;
        RECT  17.075 0.395 17.235 0.945 ;
        RECT  17.075 1.805 17.235 2.440 ;
        RECT  15.840 0.395 17.075 0.555 ;
        RECT  16.465 2.130 17.075 2.290 ;
        RECT  16.735 0.735 16.895 1.465 ;
        RECT  15.785 0.735 16.735 0.895 ;
        RECT  16.305 2.130 16.465 2.390 ;
        RECT  16.125 1.080 16.225 1.340 ;
        RECT  15.965 1.080 16.125 2.470 ;
        RECT  14.855 2.310 15.965 2.470 ;
        RECT  15.680 0.340 15.840 0.555 ;
        RECT  15.625 0.735 15.785 2.040 ;
        RECT  15.105 0.340 15.680 0.500 ;
        RECT  15.285 0.685 15.445 2.020 ;
        RECT  14.975 1.860 15.285 2.020 ;
        RECT  14.945 0.340 15.105 1.255 ;
        RECT  14.515 1.435 14.985 1.595 ;
        RECT  14.425 1.095 14.945 1.255 ;
        RECT  14.695 2.310 14.855 2.560 ;
        RECT  13.280 2.400 14.695 2.560 ;
        RECT  14.355 1.435 14.515 2.220 ;
        RECT  14.265 0.310 14.425 1.255 ;
        RECT  13.615 2.060 14.355 2.220 ;
        RECT  13.175 0.310 14.265 0.470 ;
        RECT  14.085 1.720 14.175 1.880 ;
        RECT  13.925 0.685 14.085 1.880 ;
        RECT  13.770 1.100 13.925 1.360 ;
        RECT  13.895 1.720 13.925 1.880 ;
        RECT  13.590 1.645 13.615 2.220 ;
        RECT  13.455 0.655 13.590 2.220 ;
        RECT  13.430 0.655 13.455 1.805 ;
        RECT  13.355 0.655 13.430 0.915 ;
        RECT  12.625 1.645 13.430 1.805 ;
        RECT  13.120 2.280 13.280 2.560 ;
        RECT  12.155 1.165 13.250 1.325 ;
        RECT  13.015 0.310 13.175 0.985 ;
        RECT  12.405 2.280 13.120 2.440 ;
        RECT  12.495 0.825 13.015 0.985 ;
        RECT  12.335 0.310 12.495 0.985 ;
        RECT  12.145 2.280 12.405 2.475 ;
        RECT  11.475 0.310 12.335 0.470 ;
        RECT  11.995 0.650 12.155 1.945 ;
        RECT  11.815 2.280 12.145 2.440 ;
        RECT  11.655 0.650 11.995 0.810 ;
        RECT  11.655 0.995 11.815 2.440 ;
        RECT  9.525 1.615 11.655 1.775 ;
        RECT  11.315 0.310 11.475 1.435 ;
        RECT  9.865 1.275 11.315 1.435 ;
        RECT  10.775 1.955 10.935 2.485 ;
        RECT  9.865 1.955 10.775 2.115 ;
        RECT  9.705 0.440 9.865 1.435 ;
        RECT  9.705 1.955 9.865 2.375 ;
        RECT  8.760 0.440 9.705 0.600 ;
        RECT  9.185 2.215 9.705 2.375 ;
        RECT  9.365 0.815 9.525 2.035 ;
        RECT  8.725 0.815 9.365 0.975 ;
        RECT  9.025 1.905 9.185 2.375 ;
        RECT  8.505 1.905 9.025 2.065 ;
        RECT  8.600 0.390 8.760 0.600 ;
        RECT  6.930 0.390 8.600 0.550 ;
        RECT  8.345 1.905 8.505 2.560 ;
        RECT  8.260 0.735 8.420 1.710 ;
        RECT  5.860 2.400 8.345 2.560 ;
        RECT  8.165 1.550 8.260 1.710 ;
        RECT  8.005 1.550 8.165 2.220 ;
        RECT  7.920 0.990 8.080 1.370 ;
        RECT  6.200 2.060 8.005 2.220 ;
        RECT  7.270 0.990 7.920 1.150 ;
        RECT  7.110 0.735 7.270 1.150 ;
        RECT  6.980 1.720 7.150 1.880 ;
        RECT  6.980 0.990 7.110 1.150 ;
        RECT  6.820 0.990 6.980 1.880 ;
        RECT  6.770 0.390 6.930 0.810 ;
        RECT  6.720 1.220 6.820 1.480 ;
        RECT  6.540 0.650 6.770 0.810 ;
        RECT  6.540 1.720 6.640 1.880 ;
        RECT  6.200 0.310 6.590 0.470 ;
        RECT  6.380 0.650 6.540 1.880 ;
        RECT  6.040 0.310 6.200 2.220 ;
        RECT  5.700 0.430 5.860 1.870 ;
        RECT  5.700 2.060 5.860 2.560 ;
        RECT  3.825 0.430 5.700 0.590 ;
        RECT  5.600 1.710 5.700 1.870 ;
        RECT  3.180 2.060 5.700 2.220 ;
        RECT  1.575 2.400 5.515 2.560 ;
        RECT  5.160 0.770 5.350 1.870 ;
        RECT  5.080 0.770 5.160 0.930 ;
        RECT  5.030 1.710 5.160 1.870 ;
        RECT  4.165 0.770 4.345 0.930 ;
        RECT  4.165 1.720 4.255 1.880 ;
        RECT  4.005 0.770 4.165 1.880 ;
        RECT  3.965 1.720 4.005 1.880 ;
        RECT  3.745 0.430 3.825 1.540 ;
        RECT  3.665 0.430 3.745 1.880 ;
        RECT  3.625 0.495 3.665 0.755 ;
        RECT  3.585 1.380 3.665 1.880 ;
        RECT  3.485 1.720 3.585 1.880 ;
        RECT  3.445 0.875 3.485 1.135 ;
        RECT  3.285 0.310 3.445 1.135 ;
        RECT  1.965 0.310 3.285 0.470 ;
        RECT  3.105 1.955 3.180 2.220 ;
        RECT  2.945 0.650 3.105 2.220 ;
        RECT  2.595 1.620 2.755 2.220 ;
        RECT  1.905 2.060 2.595 2.220 ;
        RECT  2.415 0.700 2.585 0.860 ;
        RECT  2.255 0.700 2.415 1.880 ;
        RECT  2.155 1.720 2.255 1.880 ;
        RECT  1.805 0.310 1.965 0.995 ;
        RECT  1.745 1.900 1.905 2.220 ;
        RECT  1.120 0.835 1.805 0.995 ;
        RECT  1.120 1.900 1.745 2.060 ;
        RECT  1.415 2.280 1.575 2.560 ;
        RECT  0.385 2.280 1.415 2.440 ;
        RECT  0.960 0.835 1.120 2.060 ;
        RECT  0.465 1.720 0.960 1.880 ;
        RECT  0.620 0.590 0.780 1.525 ;
        RECT  0.285 1.365 0.620 1.525 ;
        RECT  0.285 2.280 0.385 2.465 ;
        RECT  0.125 1.365 0.285 2.465 ;
    END
END SEDFFTRX1MTH

MACRO SEDFFTRX2MTH
    CLASS CORE ;
    FOREIGN SEDFFTRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.860 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 1.175 2.075 1.540 ;
        RECT  1.720 1.175 1.975 1.720 ;
        END
        AntennaGateArea 0.052 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 1.175 1.540 1.720 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.790 0.440 1.170 ;
        END
        AntennaGateArea 0.0624 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.730 0.405 17.940 2.080 ;
        RECT  17.545 0.405 17.730 0.565 ;
        RECT  17.585 1.820 17.730 2.080 ;
        END
        AntennaDiffArea 0.502 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.600 0.425 18.760 2.325 ;
        RECT  18.475 0.425 18.600 1.025 ;
        RECT  18.525 1.670 18.600 2.325 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.430 1.330 7.730 1.820 ;
        RECT  7.160 1.330 7.430 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 1.190 4.975 1.450 ;
        RECT  4.520 1.190 4.910 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 1.205 9.185 1.725 ;
        END
        AntennaGateArea 0.0923 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.245 -0.130 18.860 0.130 ;
        RECT  17.085 -0.130 17.245 0.380 ;
        RECT  14.765 -0.130 17.085 0.130 ;
        RECT  14.605 -0.130 14.765 0.915 ;
        RECT  12.835 -0.130 14.605 0.130 ;
        RECT  12.675 -0.130 12.835 0.645 ;
        RECT  11.135 -0.130 12.675 0.130 ;
        RECT  10.915 -0.130 11.135 1.025 ;
        RECT  10.185 -0.130 10.915 0.130 ;
        RECT  9.245 -0.130 10.185 0.250 ;
        RECT  5.110 -0.130 9.245 0.130 ;
        RECT  4.510 -0.130 5.110 0.250 ;
        RECT  1.570 -0.130 4.510 0.130 ;
        RECT  1.070 -0.130 1.570 0.300 ;
        RECT  0.725 -0.130 1.070 0.130 ;
        RECT  0.125 -0.130 0.725 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.225 2.740 18.860 3.000 ;
        RECT  16.625 2.620 17.225 3.000 ;
        RECT  12.935 2.740 16.625 3.000 ;
        RECT  12.675 2.620 12.935 3.000 ;
        RECT  10.645 2.740 12.675 3.000 ;
        RECT  10.045 2.295 10.645 3.000 ;
        RECT  8.845 2.740 10.045 3.000 ;
        RECT  8.685 2.245 8.845 3.000 ;
        RECT  1.245 2.740 8.685 3.000 ;
        RECT  0.985 2.620 1.245 3.000 ;
        RECT  0.000 2.740 0.985 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.280 1.205 18.405 1.465 ;
        RECT  18.120 1.205 18.280 2.440 ;
        RECT  17.235 2.280 18.120 2.440 ;
        RECT  17.295 0.815 17.405 1.965 ;
        RECT  17.245 0.670 17.295 1.965 ;
        RECT  17.115 0.670 17.245 1.025 ;
        RECT  17.235 1.805 17.245 1.965 ;
        RECT  17.075 1.805 17.235 2.440 ;
        RECT  16.905 0.670 17.115 0.830 ;
        RECT  16.465 2.130 17.075 2.290 ;
        RECT  16.845 1.310 17.065 1.570 ;
        RECT  16.745 0.340 16.905 0.830 ;
        RECT  16.565 1.310 16.845 1.470 ;
        RECT  15.105 0.340 16.745 0.500 ;
        RECT  16.405 0.705 16.565 1.470 ;
        RECT  16.305 2.130 16.465 2.390 ;
        RECT  15.785 0.705 16.405 0.865 ;
        RECT  16.125 1.055 16.225 1.340 ;
        RECT  15.965 1.055 16.125 2.560 ;
        RECT  13.280 2.400 15.965 2.560 ;
        RECT  15.625 0.705 15.785 2.040 ;
        RECT  15.285 0.685 15.445 2.020 ;
        RECT  14.975 1.860 15.285 2.020 ;
        RECT  14.945 0.340 15.105 1.255 ;
        RECT  14.515 1.435 14.985 1.595 ;
        RECT  14.425 1.095 14.945 1.255 ;
        RECT  14.355 1.435 14.515 2.220 ;
        RECT  14.265 0.310 14.425 1.255 ;
        RECT  13.615 2.060 14.355 2.220 ;
        RECT  13.175 0.310 14.265 0.470 ;
        RECT  14.085 1.720 14.175 1.880 ;
        RECT  13.915 0.685 14.085 1.880 ;
        RECT  13.770 1.100 13.915 1.360 ;
        RECT  13.590 1.645 13.615 2.220 ;
        RECT  13.455 0.655 13.590 2.220 ;
        RECT  13.430 0.655 13.455 1.805 ;
        RECT  13.355 0.655 13.430 0.915 ;
        RECT  12.625 1.645 13.430 1.805 ;
        RECT  13.120 2.280 13.280 2.560 ;
        RECT  12.155 1.165 13.250 1.325 ;
        RECT  13.015 0.310 13.175 0.985 ;
        RECT  12.405 2.280 13.120 2.440 ;
        RECT  12.495 0.825 13.015 0.985 ;
        RECT  12.335 0.310 12.495 0.985 ;
        RECT  12.145 2.280 12.405 2.475 ;
        RECT  11.475 0.310 12.335 0.470 ;
        RECT  11.995 0.650 12.155 1.945 ;
        RECT  11.815 2.280 12.145 2.440 ;
        RECT  11.655 0.650 11.995 0.810 ;
        RECT  11.655 0.995 11.815 2.440 ;
        RECT  9.525 1.615 11.655 1.775 ;
        RECT  11.315 0.310 11.475 1.435 ;
        RECT  11.195 1.955 11.355 2.485 ;
        RECT  9.865 1.275 11.315 1.435 ;
        RECT  9.865 1.955 11.195 2.115 ;
        RECT  9.705 0.440 9.865 1.435 ;
        RECT  9.705 1.955 9.865 2.375 ;
        RECT  8.760 0.440 9.705 0.600 ;
        RECT  9.185 2.215 9.705 2.375 ;
        RECT  9.365 0.815 9.525 2.035 ;
        RECT  8.725 0.815 9.365 0.975 ;
        RECT  9.025 1.905 9.185 2.375 ;
        RECT  8.505 1.905 9.025 2.065 ;
        RECT  8.600 0.395 8.760 0.600 ;
        RECT  6.930 0.395 8.600 0.555 ;
        RECT  8.345 1.905 8.505 2.560 ;
        RECT  8.260 0.735 8.420 1.710 ;
        RECT  5.860 2.400 8.345 2.560 ;
        RECT  8.165 1.550 8.260 1.710 ;
        RECT  8.005 1.550 8.165 2.220 ;
        RECT  7.920 0.990 8.080 1.370 ;
        RECT  6.200 2.060 8.005 2.220 ;
        RECT  7.270 0.990 7.920 1.150 ;
        RECT  7.110 0.735 7.270 1.150 ;
        RECT  6.980 1.720 7.150 1.880 ;
        RECT  6.980 0.990 7.110 1.150 ;
        RECT  6.820 0.990 6.980 1.880 ;
        RECT  6.770 0.395 6.930 0.810 ;
        RECT  6.720 1.220 6.820 1.480 ;
        RECT  6.540 0.650 6.770 0.810 ;
        RECT  6.540 1.720 6.640 1.880 ;
        RECT  6.200 0.310 6.590 0.470 ;
        RECT  6.380 0.650 6.540 1.880 ;
        RECT  6.040 0.310 6.200 2.220 ;
        RECT  5.700 0.430 5.860 1.870 ;
        RECT  5.700 2.060 5.860 2.560 ;
        RECT  3.825 0.430 5.700 0.590 ;
        RECT  5.600 1.710 5.700 1.870 ;
        RECT  3.170 2.060 5.700 2.220 ;
        RECT  1.575 2.400 5.515 2.560 ;
        RECT  5.155 0.770 5.345 1.870 ;
        RECT  5.080 0.770 5.155 0.930 ;
        RECT  5.030 1.710 5.155 1.870 ;
        RECT  4.165 0.770 4.345 0.930 ;
        RECT  4.165 1.720 4.255 1.880 ;
        RECT  4.005 0.770 4.165 1.880 ;
        RECT  3.965 1.720 4.005 1.880 ;
        RECT  3.745 0.430 3.825 1.540 ;
        RECT  3.665 0.430 3.745 1.880 ;
        RECT  3.625 0.505 3.665 0.765 ;
        RECT  3.585 1.380 3.665 1.880 ;
        RECT  3.485 1.720 3.585 1.880 ;
        RECT  3.445 0.875 3.475 1.135 ;
        RECT  3.285 0.310 3.445 1.135 ;
        RECT  1.930 0.310 3.285 0.470 ;
        RECT  3.105 1.955 3.170 2.220 ;
        RECT  2.945 0.650 3.105 2.220 ;
        RECT  2.595 1.650 2.755 2.220 ;
        RECT  1.905 2.060 2.595 2.220 ;
        RECT  2.415 0.700 2.550 0.860 ;
        RECT  2.255 0.700 2.415 1.880 ;
        RECT  2.155 1.720 2.255 1.880 ;
        RECT  1.770 0.310 1.930 0.995 ;
        RECT  1.745 1.900 1.905 2.220 ;
        RECT  1.120 0.835 1.770 0.995 ;
        RECT  1.120 1.900 1.745 2.060 ;
        RECT  1.415 2.280 1.575 2.560 ;
        RECT  0.385 2.280 1.415 2.440 ;
        RECT  0.960 0.835 1.120 2.060 ;
        RECT  0.465 1.720 0.960 1.880 ;
        RECT  0.620 0.590 0.780 1.525 ;
        RECT  0.285 1.365 0.620 1.525 ;
        RECT  0.285 2.280 0.385 2.465 ;
        RECT  0.125 1.365 0.285 2.465 ;
    END
END SEDFFTRX2MTH

MACRO SEDFFTRX4MTH
    CLASS CORE ;
    FOREIGN SEDFFTRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.090 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.960 1.200 2.075 1.460 ;
        RECT  1.720 1.175 1.960 1.720 ;
        END
        AntennaGateArea 0.052 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.300 1.175 1.540 1.720 ;
        END
        AntennaGateArea 0.1157 ;
    END SE
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.790 0.440 1.170 ;
        END
        AntennaGateArea 0.0624 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.115 0.425 18.375 1.895 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.405 1.290 19.705 1.580 ;
        RECT  19.405 0.425 19.455 1.025 ;
        RECT  19.245 0.425 19.405 2.425 ;
        RECT  19.195 0.425 19.245 1.025 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.425 1.330 7.730 1.750 ;
        RECT  7.160 1.330 7.425 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.910 1.190 4.970 1.450 ;
        RECT  4.520 1.190 4.910 1.540 ;
        END
        AntennaGateArea 0.0533 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.710 1.205 9.185 1.725 ;
        END
        AntennaGateArea 0.1053 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.965 -0.130 20.090 0.130 ;
        RECT  19.705 -0.130 19.965 1.025 ;
        RECT  18.945 -0.130 19.705 0.130 ;
        RECT  18.685 -0.130 18.945 1.025 ;
        RECT  17.865 -0.130 18.685 0.130 ;
        RECT  17.605 -0.130 17.865 0.660 ;
        RECT  14.765 -0.130 17.605 0.130 ;
        RECT  14.605 -0.130 14.765 0.915 ;
        RECT  12.835 -0.130 14.605 0.130 ;
        RECT  12.675 -0.130 12.835 0.645 ;
        RECT  11.135 -0.130 12.675 0.130 ;
        RECT  10.915 -0.130 11.135 1.025 ;
        RECT  10.185 -0.130 10.915 0.130 ;
        RECT  9.245 -0.130 10.185 0.250 ;
        RECT  5.110 -0.130 9.245 0.130 ;
        RECT  4.510 -0.130 5.110 0.250 ;
        RECT  1.450 -0.130 4.510 0.130 ;
        RECT  1.190 -0.130 1.450 0.305 ;
        RECT  0.725 -0.130 1.190 0.130 ;
        RECT  0.125 -0.130 0.725 0.250 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.915 2.740 20.090 3.000 ;
        RECT  19.755 1.825 19.915 3.000 ;
        RECT  18.915 2.740 19.755 3.000 ;
        RECT  18.655 2.420 18.915 3.000 ;
        RECT  17.835 2.740 18.655 3.000 ;
        RECT  17.575 2.620 17.835 3.000 ;
        RECT  16.785 2.740 17.575 3.000 ;
        RECT  16.525 2.620 16.785 3.000 ;
        RECT  12.935 2.740 16.525 3.000 ;
        RECT  12.675 2.620 12.935 3.000 ;
        RECT  10.645 2.740 12.675 3.000 ;
        RECT  10.045 2.295 10.645 3.000 ;
        RECT  8.845 2.740 10.045 3.000 ;
        RECT  8.685 2.245 8.845 3.000 ;
        RECT  1.245 2.740 8.685 3.000 ;
        RECT  0.985 2.620 1.245 3.000 ;
        RECT  0.000 2.740 0.985 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  18.905 1.205 19.065 2.235 ;
        RECT  17.815 2.075 18.905 2.235 ;
        RECT  17.655 0.870 17.815 2.235 ;
        RECT  17.295 0.870 17.655 1.030 ;
        RECT  17.285 2.075 17.655 2.235 ;
        RECT  16.895 1.240 17.465 1.500 ;
        RECT  17.135 0.310 17.295 1.030 ;
        RECT  17.115 1.900 17.285 2.235 ;
        RECT  15.105 0.310 17.135 0.470 ;
        RECT  16.470 2.035 17.115 2.235 ;
        RECT  16.735 0.665 16.895 1.500 ;
        RECT  15.785 0.665 16.735 0.825 ;
        RECT  16.310 2.035 16.470 2.320 ;
        RECT  16.125 1.035 16.265 1.195 ;
        RECT  15.965 1.035 16.125 2.560 ;
        RECT  13.280 2.400 15.965 2.560 ;
        RECT  15.625 0.665 15.785 2.040 ;
        RECT  15.285 0.685 15.445 2.020 ;
        RECT  14.975 1.860 15.285 2.020 ;
        RECT  14.945 0.310 15.105 1.255 ;
        RECT  14.515 1.435 14.985 1.595 ;
        RECT  14.425 1.095 14.945 1.255 ;
        RECT  14.355 1.435 14.515 2.220 ;
        RECT  14.265 0.310 14.425 1.255 ;
        RECT  13.615 2.060 14.355 2.220 ;
        RECT  13.175 0.310 14.265 0.470 ;
        RECT  14.085 1.720 14.175 1.880 ;
        RECT  13.915 0.685 14.085 1.880 ;
        RECT  13.770 1.100 13.915 1.360 ;
        RECT  13.590 1.645 13.615 2.220 ;
        RECT  13.455 0.670 13.590 2.220 ;
        RECT  13.430 0.670 13.455 1.805 ;
        RECT  13.355 0.670 13.430 0.930 ;
        RECT  12.625 1.645 13.430 1.805 ;
        RECT  13.120 2.280 13.280 2.560 ;
        RECT  12.155 1.165 13.250 1.325 ;
        RECT  13.015 0.310 13.175 0.985 ;
        RECT  12.405 2.280 13.120 2.440 ;
        RECT  12.495 0.825 13.015 0.985 ;
        RECT  12.335 0.310 12.495 0.985 ;
        RECT  12.145 2.280 12.405 2.475 ;
        RECT  11.475 0.310 12.335 0.470 ;
        RECT  11.995 0.650 12.155 1.945 ;
        RECT  11.815 2.280 12.145 2.440 ;
        RECT  11.655 0.650 11.995 0.810 ;
        RECT  11.655 0.995 11.815 2.440 ;
        RECT  9.525 1.615 11.655 1.775 ;
        RECT  11.315 0.310 11.475 1.435 ;
        RECT  11.195 1.955 11.355 2.485 ;
        RECT  9.865 1.275 11.315 1.435 ;
        RECT  9.865 1.955 11.195 2.115 ;
        RECT  9.705 0.440 9.865 1.435 ;
        RECT  9.705 1.955 9.865 2.375 ;
        RECT  8.760 0.440 9.705 0.600 ;
        RECT  9.185 2.215 9.705 2.375 ;
        RECT  9.365 0.815 9.525 2.035 ;
        RECT  8.725 0.815 9.365 0.975 ;
        RECT  9.025 1.905 9.185 2.375 ;
        RECT  8.505 1.905 9.025 2.065 ;
        RECT  8.600 0.395 8.760 0.600 ;
        RECT  6.930 0.395 8.600 0.555 ;
        RECT  8.345 1.905 8.505 2.560 ;
        RECT  8.260 0.735 8.420 1.710 ;
        RECT  5.860 2.400 8.345 2.560 ;
        RECT  8.165 1.550 8.260 1.710 ;
        RECT  8.005 1.550 8.165 2.220 ;
        RECT  7.920 0.990 8.080 1.370 ;
        RECT  6.200 2.060 8.005 2.220 ;
        RECT  7.270 0.990 7.920 1.150 ;
        RECT  7.110 0.735 7.270 1.150 ;
        RECT  6.980 1.720 7.150 1.880 ;
        RECT  6.980 0.990 7.110 1.150 ;
        RECT  6.820 0.990 6.980 1.880 ;
        RECT  6.770 0.395 6.930 0.810 ;
        RECT  6.720 1.220 6.820 1.480 ;
        RECT  6.540 0.650 6.770 0.810 ;
        RECT  6.540 1.720 6.640 1.880 ;
        RECT  6.200 0.310 6.590 0.470 ;
        RECT  6.380 0.650 6.540 1.880 ;
        RECT  6.040 0.310 6.200 2.220 ;
        RECT  5.700 0.430 5.860 1.870 ;
        RECT  5.700 2.060 5.860 2.560 ;
        RECT  3.825 0.430 5.700 0.590 ;
        RECT  5.600 1.710 5.700 1.870 ;
        RECT  3.170 2.060 5.700 2.220 ;
        RECT  1.575 2.400 5.515 2.560 ;
        RECT  5.150 0.770 5.340 1.870 ;
        RECT  5.080 0.770 5.150 0.930 ;
        RECT  5.030 1.710 5.150 1.870 ;
        RECT  4.165 0.770 4.340 0.930 ;
        RECT  4.165 1.720 4.255 1.880 ;
        RECT  4.005 0.770 4.165 1.880 ;
        RECT  3.965 1.720 4.005 1.880 ;
        RECT  3.785 0.430 3.825 1.375 ;
        RECT  3.695 0.365 3.785 1.375 ;
        RECT  3.695 1.720 3.745 1.880 ;
        RECT  3.665 0.365 3.695 1.880 ;
        RECT  3.625 0.365 3.665 0.625 ;
        RECT  3.535 1.215 3.665 1.880 ;
        RECT  3.485 1.720 3.535 1.880 ;
        RECT  3.445 0.775 3.485 1.035 ;
        RECT  3.285 0.310 3.445 1.035 ;
        RECT  1.965 0.310 3.285 0.470 ;
        RECT  3.105 1.955 3.170 2.220 ;
        RECT  2.945 0.650 3.105 2.220 ;
        RECT  2.595 1.620 2.755 2.220 ;
        RECT  1.905 2.060 2.595 2.220 ;
        RECT  2.415 0.700 2.585 0.860 ;
        RECT  2.255 0.700 2.415 1.880 ;
        RECT  2.155 1.720 2.255 1.880 ;
        RECT  1.805 0.310 1.965 0.995 ;
        RECT  1.745 1.900 1.905 2.220 ;
        RECT  1.120 0.835 1.805 0.995 ;
        RECT  1.120 1.900 1.745 2.060 ;
        RECT  1.415 2.280 1.575 2.560 ;
        RECT  0.385 2.280 1.415 2.440 ;
        RECT  0.960 0.835 1.120 2.060 ;
        RECT  0.465 1.720 0.960 1.880 ;
        RECT  0.620 0.590 0.780 1.525 ;
        RECT  0.285 1.365 0.620 1.525 ;
        RECT  0.285 2.280 0.385 2.465 ;
        RECT  0.125 1.365 0.285 2.465 ;
    END
END SEDFFTRX4MTH

MACRO SEDFFX1MTH
    CLASS CORE ;
    FOREIGN SEDFFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.580 1.620 1.915 1.780 ;
        RECT  1.355 1.620 1.580 1.950 ;
        RECT  1.290 1.740 1.355 1.950 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.405 1.640 ;
        END
        AntennaGateArea 0.1365 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.200 1.755 12.745 2.015 ;
        RECT  12.200 0.815 12.710 1.025 ;
        RECT  11.990 0.815 12.200 2.015 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 1.290 14.250 1.580 ;
        RECT  13.950 0.760 14.225 1.925 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.195 5.015 1.540 ;
        RECT  4.610 1.195 4.820 1.580 ;
        RECT  3.700 1.380 4.610 1.540 ;
        RECT  3.540 1.380 3.700 1.725 ;
        END
        AntennaGateArea 0.1378 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.095 2.870 1.540 ;
        END
        AntennaGateArea 0.0845 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.670 1.070 9.060 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.565 -0.130 14.350 0.130 ;
        RECT  12.965 -0.130 13.565 0.250 ;
        RECT  12.600 -0.130 12.965 0.130 ;
        RECT  12.000 -0.130 12.600 0.250 ;
        RECT  10.580 -0.130 12.000 0.130 ;
        RECT  10.320 -0.130 10.580 0.300 ;
        RECT  7.545 -0.130 10.320 0.130 ;
        RECT  7.385 -0.130 7.545 0.300 ;
        RECT  5.270 -0.130 7.385 0.130 ;
        RECT  5.010 -0.130 5.270 0.250 ;
        RECT  1.910 -0.130 5.010 0.130 ;
        RECT  1.650 -0.130 1.910 0.575 ;
        RECT  0.725 -0.130 1.650 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  14.005 2.740 14.350 3.000 ;
        RECT  13.405 2.565 14.005 3.000 ;
        RECT  12.980 2.740 13.405 3.000 ;
        RECT  12.380 2.565 12.980 3.000 ;
        RECT  1.795 2.740 12.380 3.000 ;
        RECT  1.535 2.570 1.795 3.000 ;
        RECT  0.385 2.740 1.535 3.000 ;
        RECT  0.125 2.470 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.720 1.230 13.770 1.490 ;
        RECT  13.510 0.430 13.720 1.490 ;
        RECT  11.815 0.430 13.510 0.590 ;
        RECT  13.205 0.815 13.285 0.975 ;
        RECT  13.045 0.815 13.205 2.360 ;
        RECT  12.960 0.815 13.045 0.975 ;
        RECT  12.380 1.260 13.045 1.520 ;
        RECT  12.150 2.200 13.045 2.360 ;
        RECT  11.990 2.200 12.150 2.560 ;
        RECT  4.520 2.400 11.990 2.560 ;
        RECT  11.810 0.355 11.815 0.590 ;
        RECT  11.650 0.355 11.810 2.220 ;
        RECT  10.950 0.355 11.650 0.515 ;
        RECT  11.195 1.960 11.650 2.220 ;
        RECT  11.285 0.840 11.470 1.100 ;
        RECT  11.125 0.695 11.285 1.780 ;
        RECT  10.140 0.695 11.125 0.855 ;
        RECT  10.985 1.620 11.125 1.780 ;
        RECT  10.825 1.620 10.985 2.220 ;
        RECT  10.645 1.155 10.945 1.415 ;
        RECT  6.515 2.060 10.825 2.220 ;
        RECT  10.485 1.035 10.645 1.880 ;
        RECT  9.800 1.035 10.485 1.195 ;
        RECT  9.675 1.720 10.485 1.880 ;
        RECT  9.420 1.380 10.305 1.540 ;
        RECT  9.980 0.310 10.140 0.855 ;
        RECT  9.290 0.310 9.980 0.470 ;
        RECT  9.640 0.680 9.800 1.195 ;
        RECT  9.540 0.680 9.640 0.890 ;
        RECT  8.830 0.730 9.540 0.890 ;
        RECT  9.260 1.380 9.420 1.880 ;
        RECT  9.030 0.310 9.290 0.520 ;
        RECT  8.490 1.720 9.260 1.880 ;
        RECT  8.670 0.325 8.830 0.890 ;
        RECT  7.885 0.325 8.670 0.485 ;
        RECT  8.330 0.690 8.490 1.880 ;
        RECT  8.065 0.690 8.330 0.850 ;
        RECT  7.600 1.720 8.330 1.880 ;
        RECT  7.870 1.030 8.030 1.490 ;
        RECT  7.725 0.325 7.885 0.650 ;
        RECT  6.855 1.030 7.870 1.190 ;
        RECT  7.195 0.490 7.725 0.650 ;
        RECT  7.440 1.370 7.600 1.880 ;
        RECT  7.340 1.370 7.440 1.575 ;
        RECT  7.035 0.325 7.195 0.650 ;
        RECT  6.780 0.325 7.035 0.485 ;
        RECT  6.695 0.695 6.855 1.880 ;
        RECT  6.550 0.695 6.695 0.855 ;
        RECT  6.370 1.115 6.515 2.220 ;
        RECT  6.355 0.720 6.370 2.220 ;
        RECT  6.210 0.720 6.355 1.275 ;
        RECT  6.055 0.355 6.240 0.515 ;
        RECT  6.015 1.810 6.175 2.220 ;
        RECT  5.895 0.355 6.055 0.590 ;
        RECT  4.410 2.060 6.015 2.220 ;
        RECT  4.755 0.430 5.895 0.590 ;
        RECT  5.570 0.790 5.730 1.880 ;
        RECT  5.450 0.790 5.570 1.020 ;
        RECT  4.950 1.720 5.570 1.880 ;
        RECT  4.430 0.790 5.450 0.950 ;
        RECT  4.495 0.355 4.755 0.590 ;
        RECT  4.090 0.430 4.495 0.590 ;
        RECT  4.270 0.790 4.430 1.195 ;
        RECT  4.200 2.015 4.410 2.220 ;
        RECT  3.210 1.035 4.270 1.195 ;
        RECT  3.030 2.015 4.200 2.175 ;
        RECT  3.930 0.430 4.090 0.855 ;
        RECT  2.560 0.695 3.930 0.855 ;
        RECT  2.295 0.355 3.750 0.515 ;
        RECT  3.245 2.355 3.505 2.560 ;
        RECT  2.165 2.400 3.245 2.560 ;
        RECT  3.050 1.035 3.210 1.835 ;
        RECT  2.870 2.015 3.030 2.220 ;
        RECT  2.345 2.060 2.870 2.220 ;
        RECT  2.280 1.690 2.395 1.850 ;
        RECT  2.135 0.355 2.295 0.915 ;
        RECT  2.120 1.120 2.280 1.850 ;
        RECT  2.005 2.180 2.165 2.560 ;
        RECT  1.340 0.755 2.135 0.915 ;
        RECT  0.830 1.120 2.120 1.280 ;
        RECT  1.225 2.180 2.005 2.340 ;
        RECT  1.095 0.645 1.340 0.915 ;
        RECT  0.965 2.180 1.225 2.465 ;
        RECT  0.825 0.815 0.830 1.280 ;
        RECT  0.665 0.815 0.825 2.030 ;
        RECT  0.570 0.815 0.665 0.975 ;
        RECT  0.565 1.765 0.665 2.030 ;
    END
END SEDFFX1MTH

MACRO SEDFFX2MTH
    CLASS CORE ;
    FOREIGN SEDFFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.350 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.285 1.620 1.875 1.950 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.075 0.445 1.620 ;
        END
        AntennaGateArea 0.1365 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.225 1.290 14.250 1.580 ;
        RECT  13.965 0.400 14.225 2.355 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.315 0.880 13.430 1.170 ;
        RECT  13.055 0.765 13.315 1.925 ;
        END
        AntennaDiffArea 0.438 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.875 1.195 5.300 1.540 ;
        RECT  4.610 1.195 4.875 1.580 ;
        RECT  3.700 1.380 4.610 1.540 ;
        RECT  3.540 1.380 3.700 1.835 ;
        END
        AntennaGateArea 0.1378 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.095 2.870 1.540 ;
        END
        AntennaGateArea 0.0845 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.670 1.090 9.060 1.540 ;
        END
        AntennaGateArea 0.0884 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.690 -0.130 14.350 0.130 ;
        RECT  13.430 -0.130 13.690 0.535 ;
        RECT  12.655 -0.130 13.430 0.130 ;
        RECT  12.055 -0.130 12.655 0.250 ;
        RECT  10.480 -0.130 12.055 0.130 ;
        RECT  10.320 -0.130 10.480 0.300 ;
        RECT  7.570 -0.130 10.320 0.130 ;
        RECT  7.410 -0.130 7.570 0.300 ;
        RECT  5.260 -0.130 7.410 0.130 ;
        RECT  5.000 -0.130 5.260 0.250 ;
        RECT  1.910 -0.130 5.000 0.130 ;
        RECT  1.650 -0.130 1.910 0.575 ;
        RECT  0.725 -0.130 1.650 0.130 ;
        RECT  0.125 -0.130 0.725 0.365 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.745 2.740 14.350 3.000 ;
        RECT  12.145 2.470 12.745 3.000 ;
        RECT  1.795 2.740 12.145 3.000 ;
        RECT  1.535 2.570 1.795 3.000 ;
        RECT  0.385 2.740 1.535 3.000 ;
        RECT  0.125 2.470 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.615 1.270 13.775 2.265 ;
        RECT  12.295 2.105 13.615 2.265 ;
        RECT  12.760 1.200 12.860 1.460 ;
        RECT  12.600 0.430 12.760 1.460 ;
        RECT  11.815 0.430 12.600 0.595 ;
        RECT  12.295 0.815 12.370 0.975 ;
        RECT  12.135 0.815 12.295 2.265 ;
        RECT  12.055 0.815 12.135 0.975 ;
        RECT  11.995 1.310 12.135 1.570 ;
        RECT  11.965 2.105 12.135 2.265 ;
        RECT  11.805 2.105 11.965 2.560 ;
        RECT  11.655 0.355 11.815 1.790 ;
        RECT  4.520 2.400 11.805 2.560 ;
        RECT  10.950 0.355 11.655 0.515 ;
        RECT  11.625 1.630 11.655 1.790 ;
        RECT  11.465 1.630 11.625 2.220 ;
        RECT  11.285 0.845 11.470 1.105 ;
        RECT  11.165 2.060 11.465 2.220 ;
        RECT  11.125 0.695 11.285 1.850 ;
        RECT  10.140 0.695 11.125 0.855 ;
        RECT  10.985 1.690 11.125 1.850 ;
        RECT  10.825 1.690 10.985 2.220 ;
        RECT  10.645 1.155 10.945 1.415 ;
        RECT  6.515 2.060 10.825 2.220 ;
        RECT  10.485 1.035 10.645 1.880 ;
        RECT  9.800 1.035 10.485 1.195 ;
        RECT  9.675 1.720 10.485 1.880 ;
        RECT  9.420 1.380 10.305 1.540 ;
        RECT  9.980 0.310 10.140 0.855 ;
        RECT  9.290 0.310 9.980 0.470 ;
        RECT  9.640 0.655 9.800 1.195 ;
        RECT  9.540 0.655 9.640 0.860 ;
        RECT  8.830 0.700 9.540 0.860 ;
        RECT  9.260 1.380 9.420 1.880 ;
        RECT  9.030 0.310 9.290 0.520 ;
        RECT  8.490 1.720 9.260 1.880 ;
        RECT  8.670 0.325 8.830 0.860 ;
        RECT  7.910 0.325 8.670 0.485 ;
        RECT  8.330 0.695 8.490 1.880 ;
        RECT  8.090 0.695 8.330 0.855 ;
        RECT  7.600 1.720 8.330 1.880 ;
        RECT  7.870 1.030 8.030 1.490 ;
        RECT  7.750 0.325 7.910 0.735 ;
        RECT  6.885 1.030 7.870 1.190 ;
        RECT  7.230 0.575 7.750 0.735 ;
        RECT  7.440 1.415 7.600 1.880 ;
        RECT  7.340 1.415 7.440 1.575 ;
        RECT  7.070 0.325 7.230 0.735 ;
        RECT  6.860 0.325 7.070 0.485 ;
        RECT  6.855 0.695 6.885 1.190 ;
        RECT  6.695 0.695 6.855 1.880 ;
        RECT  6.625 0.695 6.695 0.855 ;
        RECT  6.435 1.115 6.515 2.220 ;
        RECT  6.355 0.820 6.435 2.220 ;
        RECT  6.275 0.820 6.355 1.275 ;
        RECT  6.175 0.820 6.275 0.980 ;
        RECT  4.750 0.430 6.250 0.590 ;
        RECT  6.015 1.780 6.175 2.220 ;
        RECT  4.360 2.060 6.015 2.220 ;
        RECT  5.580 0.770 5.740 1.880 ;
        RECT  5.460 0.770 5.580 1.000 ;
        RECT  5.020 1.720 5.580 1.880 ;
        RECT  4.430 0.770 5.460 0.930 ;
        RECT  4.490 0.355 4.750 0.590 ;
        RECT  4.090 0.430 4.490 0.590 ;
        RECT  4.270 0.770 4.430 1.200 ;
        RECT  4.150 2.015 4.360 2.220 ;
        RECT  3.260 1.040 4.270 1.200 ;
        RECT  3.030 2.015 4.150 2.175 ;
        RECT  3.930 0.430 4.090 0.855 ;
        RECT  2.560 0.695 3.930 0.855 ;
        RECT  2.295 0.355 3.750 0.515 ;
        RECT  3.245 2.355 3.505 2.560 ;
        RECT  3.100 1.040 3.260 1.835 ;
        RECT  2.165 2.400 3.245 2.560 ;
        RECT  2.995 1.675 3.100 1.835 ;
        RECT  2.870 2.015 3.030 2.220 ;
        RECT  2.345 2.060 2.870 2.220 ;
        RECT  2.245 1.670 2.360 1.830 ;
        RECT  2.135 0.355 2.295 0.915 ;
        RECT  2.085 1.120 2.245 1.830 ;
        RECT  2.005 2.180 2.165 2.560 ;
        RECT  1.290 0.755 2.135 0.915 ;
        RECT  0.825 1.120 2.085 1.280 ;
        RECT  1.225 2.180 2.005 2.340 ;
        RECT  1.130 0.600 1.290 0.915 ;
        RECT  0.965 2.180 1.225 2.465 ;
        RECT  0.665 0.750 0.825 1.980 ;
        RECT  0.565 0.750 0.665 0.910 ;
        RECT  0.565 1.820 0.665 1.980 ;
    END
END SEDFFX2MTH

MACRO SEDFFX4MTH
    CLASS CORE ;
    FOREIGN SEDFFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.290 1.620 1.910 1.950 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.185 0.485 1.580 ;
        END
        AntennaGateArea 0.1378 ;
    END SE
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.700 0.425 14.940 2.300 ;
        RECT  14.665 0.425 14.700 1.025 ;
        RECT  14.680 1.700 14.700 2.300 ;
        RECT  14.450 1.700 14.680 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  13.850 0.425 13.920 1.025 ;
        RECT  13.590 0.425 13.850 1.955 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.195 5.300 1.535 ;
        RECT  4.610 1.195 4.820 1.580 ;
        RECT  3.700 1.375 4.610 1.535 ;
        RECT  3.540 1.375 3.700 1.725 ;
        END
        AntennaGateArea 0.1365 ;
    END E
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.520 1.095 2.870 1.540 ;
        END
        AntennaGateArea 0.0845 ;
    END D
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  8.670 1.070 9.060 1.540 ;
        END
        AntennaGateArea 0.1092 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.450 -0.130 15.580 0.130 ;
        RECT  15.190 -0.130 15.450 0.965 ;
        RECT  14.430 -0.130 15.190 0.130 ;
        RECT  14.170 -0.130 14.430 0.975 ;
        RECT  13.290 -0.130 14.170 0.130 ;
        RECT  12.350 -0.130 13.290 0.300 ;
        RECT  7.545 -0.130 12.350 0.130 ;
        RECT  7.385 -0.130 7.545 0.300 ;
        RECT  5.260 -0.130 7.385 0.130 ;
        RECT  5.000 -0.130 5.260 0.250 ;
        RECT  1.910 -0.130 5.000 0.130 ;
        RECT  1.650 -0.130 1.910 0.575 ;
        RECT  0.725 -0.130 1.650 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.450 2.740 15.580 3.000 ;
        RECT  15.190 1.895 15.450 3.000 ;
        RECT  14.395 2.740 15.190 3.000 ;
        RECT  14.135 2.570 14.395 3.000 ;
        RECT  13.300 2.740 14.135 3.000 ;
        RECT  12.360 2.570 13.300 3.000 ;
        RECT  4.400 2.740 12.360 3.000 ;
        RECT  3.900 2.570 4.400 3.000 ;
        RECT  1.605 2.740 3.900 3.000 ;
        RECT  1.345 2.520 1.605 3.000 ;
        RECT  0.385 2.740 1.345 3.000 ;
        RECT  0.125 1.890 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  14.360 1.200 14.520 1.465 ;
        RECT  14.190 1.300 14.360 1.465 ;
        RECT  14.030 1.300 14.190 2.295 ;
        RECT  13.410 2.135 14.030 2.295 ;
        RECT  13.250 0.705 13.410 2.295 ;
        RECT  12.680 0.705 13.250 0.940 ;
        RECT  12.230 1.900 13.250 2.160 ;
        RECT  12.455 1.120 13.060 1.465 ;
        RECT  12.160 1.120 12.455 1.280 ;
        RECT  12.130 1.460 12.230 2.160 ;
        RECT  12.000 0.310 12.160 1.280 ;
        RECT  11.970 1.460 12.130 2.560 ;
        RECT  11.160 0.310 12.000 0.470 ;
        RECT  11.790 1.120 12.000 1.280 ;
        RECT  4.615 2.400 11.970 2.560 ;
        RECT  11.630 1.120 11.790 2.220 ;
        RECT  11.395 0.650 11.655 0.855 ;
        RECT  11.280 2.060 11.630 2.220 ;
        RECT  11.390 0.695 11.395 0.855 ;
        RECT  11.230 0.695 11.390 1.750 ;
        RECT  10.300 0.695 11.230 0.855 ;
        RECT  10.985 1.590 11.230 1.750 ;
        RECT  10.900 0.310 11.160 0.515 ;
        RECT  10.825 1.590 10.985 2.220 ;
        RECT  10.645 1.095 10.910 1.355 ;
        RECT  6.515 2.060 10.825 2.220 ;
        RECT  10.485 1.035 10.645 1.880 ;
        RECT  9.800 1.035 10.485 1.195 ;
        RECT  9.675 1.720 10.485 1.880 ;
        RECT  9.420 1.380 10.305 1.540 ;
        RECT  10.140 0.310 10.300 0.855 ;
        RECT  9.290 0.310 10.140 0.470 ;
        RECT  9.640 0.650 9.800 1.195 ;
        RECT  9.540 0.650 9.640 0.860 ;
        RECT  8.830 0.700 9.540 0.860 ;
        RECT  9.260 1.380 9.420 1.880 ;
        RECT  9.030 0.310 9.290 0.520 ;
        RECT  8.490 1.720 9.260 1.880 ;
        RECT  8.670 0.325 8.830 0.860 ;
        RECT  7.890 0.325 8.670 0.485 ;
        RECT  8.330 0.665 8.490 1.880 ;
        RECT  8.090 0.665 8.330 0.825 ;
        RECT  7.600 1.720 8.330 1.880 ;
        RECT  7.870 1.030 8.030 1.490 ;
        RECT  7.730 0.325 7.890 0.645 ;
        RECT  6.855 1.030 7.870 1.190 ;
        RECT  7.200 0.485 7.730 0.645 ;
        RECT  7.440 1.415 7.600 1.880 ;
        RECT  7.340 1.415 7.440 1.575 ;
        RECT  7.040 0.325 7.200 0.645 ;
        RECT  6.780 0.325 7.040 0.485 ;
        RECT  6.695 0.695 6.855 1.880 ;
        RECT  6.550 0.695 6.695 0.855 ;
        RECT  6.370 1.115 6.515 2.220 ;
        RECT  6.355 0.800 6.370 2.220 ;
        RECT  6.110 0.800 6.355 1.275 ;
        RECT  5.980 0.355 6.240 0.605 ;
        RECT  5.945 1.960 6.175 2.220 ;
        RECT  4.750 0.445 5.980 0.605 ;
        RECT  4.410 2.060 5.945 2.220 ;
        RECT  5.570 0.785 5.730 1.880 ;
        RECT  5.450 0.785 5.570 1.015 ;
        RECT  5.020 1.720 5.570 1.880 ;
        RECT  4.430 0.785 5.450 0.945 ;
        RECT  4.490 0.355 4.750 0.605 ;
        RECT  4.090 0.445 4.490 0.605 ;
        RECT  4.270 0.785 4.430 1.195 ;
        RECT  4.150 1.960 4.410 2.220 ;
        RECT  3.260 1.035 4.270 1.195 ;
        RECT  3.030 2.015 4.150 2.175 ;
        RECT  3.930 0.445 4.090 0.855 ;
        RECT  2.560 0.695 3.930 0.855 ;
        RECT  2.295 0.355 3.750 0.515 ;
        RECT  3.245 2.355 3.505 2.560 ;
        RECT  3.100 1.035 3.260 1.835 ;
        RECT  2.155 2.400 3.245 2.560 ;
        RECT  2.995 1.675 3.100 1.835 ;
        RECT  2.870 2.015 3.030 2.220 ;
        RECT  2.345 2.060 2.870 2.220 ;
        RECT  2.280 1.690 2.395 1.850 ;
        RECT  2.135 0.355 2.295 0.915 ;
        RECT  2.120 1.120 2.280 1.850 ;
        RECT  1.995 2.180 2.155 2.560 ;
        RECT  1.340 0.755 2.135 0.915 ;
        RECT  0.825 1.120 2.120 1.280 ;
        RECT  0.955 2.180 1.995 2.340 ;
        RECT  1.080 0.600 1.340 0.915 ;
        RECT  0.825 1.735 0.965 1.895 ;
        RECT  0.695 2.180 0.955 2.485 ;
        RECT  0.665 0.815 0.825 1.895 ;
        RECT  0.565 0.815 0.665 0.975 ;
    END
END SEDFFX4MTH

MACRO SMDFFHQX1MTH
    CLASS CORE ;
    FOREIGN SMDFFHQX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.220 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.205 1.185 1.465 ;
        RECT  0.920 1.205 1.130 1.990 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 0.310 5.780 0.470 ;
        RECT  1.115 0.310 1.275 0.660 ;
        RECT  0.730 0.500 1.115 0.660 ;
        RECT  0.570 0.500 0.730 1.580 ;
        RECT  0.435 1.280 0.570 1.580 ;
        END
        AntennaGateArea 0.1469 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.985 1.230 6.245 1.420 ;
        RECT  5.640 1.260 5.985 1.420 ;
        RECT  5.430 1.260 5.640 1.580 ;
        RECT  4.810 1.260 5.430 1.420 ;
        RECT  4.650 1.160 4.810 1.420 ;
        END
        AntennaGateArea 0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.095 1.290 17.120 1.580 ;
        RECT  16.905 0.740 17.095 2.095 ;
        RECT  16.835 0.740 16.905 1.000 ;
        RECT  16.835 1.835 16.905 2.095 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 1.175 3.590 1.580 ;
        RECT  2.745 1.175 3.350 1.435 ;
        END
        AntennaGateArea 0.0611 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.375 0.470 8.510 0.770 ;
        RECT  8.215 0.470 8.375 1.250 ;
        END
        AntennaGateArea 0.0663 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.210 0.650 9.450 1.170 ;
        RECT  9.030 0.880 9.210 1.170 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.530 -0.130 17.220 0.130 ;
        RECT  16.370 -0.130 16.530 0.965 ;
        RECT  15.785 -0.130 16.370 0.300 ;
        RECT  15.565 -0.130 15.785 0.130 ;
        RECT  15.065 -0.130 15.565 0.300 ;
        RECT  13.630 -0.130 15.065 0.130 ;
        RECT  13.030 -0.130 13.630 0.355 ;
        RECT  11.190 -0.130 13.030 0.130 ;
        RECT  10.690 -0.130 11.190 0.300 ;
        RECT  9.495 -0.130 10.690 0.130 ;
        RECT  9.335 -0.130 9.495 0.300 ;
        RECT  7.190 -0.130 9.335 0.130 ;
        RECT  6.350 -0.130 7.190 0.300 ;
        RECT  0.765 -0.130 6.350 0.130 ;
        RECT  0.265 -0.130 0.765 0.300 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.425 2.740 17.220 3.000 ;
        RECT  15.585 2.400 16.425 3.000 ;
        RECT  8.050 2.740 15.585 3.000 ;
        RECT  7.450 2.620 8.050 3.000 ;
        RECT  6.490 2.740 7.450 3.000 ;
        RECT  5.550 2.620 6.490 3.000 ;
        RECT  0.755 2.740 5.550 3.000 ;
        RECT  0.255 2.570 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.030 0.600 16.190 2.110 ;
        RECT  15.800 0.600 16.030 0.760 ;
        RECT  15.945 1.575 16.030 2.110 ;
        RECT  15.455 1.575 15.945 1.735 ;
        RECT  15.650 0.940 15.810 1.235 ;
        RECT  14.915 0.940 15.650 1.100 ;
        RECT  15.295 1.460 15.455 1.735 ;
        RECT  14.925 2.365 15.025 2.525 ;
        RECT  14.765 2.060 14.925 2.525 ;
        RECT  14.755 0.575 14.915 1.855 ;
        RECT  14.385 2.060 14.765 2.220 ;
        RECT  14.745 0.575 14.755 0.735 ;
        RECT  14.565 1.695 14.755 1.855 ;
        RECT  14.485 0.545 14.745 0.735 ;
        RECT  14.385 0.915 14.575 1.145 ;
        RECT  11.670 2.400 14.405 2.560 ;
        RECT  14.315 0.915 14.385 2.220 ;
        RECT  14.225 0.985 14.315 2.220 ;
        RECT  14.135 0.545 14.235 0.705 ;
        RECT  12.010 2.060 14.225 2.220 ;
        RECT  14.045 0.545 14.135 0.760 ;
        RECT  13.975 0.545 14.045 1.860 ;
        RECT  13.885 0.600 13.975 1.860 ;
        RECT  13.225 0.600 13.885 0.760 ;
        RECT  13.785 1.700 13.885 1.860 ;
        RECT  13.605 1.030 13.705 1.290 ;
        RECT  13.445 1.030 13.605 1.810 ;
        RECT  12.885 1.650 13.445 1.810 ;
        RECT  13.065 0.600 13.225 1.265 ;
        RECT  12.725 0.645 12.885 1.810 ;
        RECT  12.355 0.645 12.725 0.805 ;
        RECT  12.355 1.650 12.725 1.810 ;
        RECT  12.010 1.010 12.535 1.270 ;
        RECT  12.195 0.545 12.355 0.805 ;
        RECT  12.195 1.620 12.355 1.880 ;
        RECT  11.850 0.620 12.010 2.220 ;
        RECT  10.975 0.620 11.850 0.780 ;
        RECT  11.510 0.990 11.670 2.560 ;
        RECT  11.180 0.990 11.510 1.150 ;
        RECT  10.980 1.960 11.510 2.120 ;
        RECT  11.170 2.300 11.330 2.560 ;
        RECT  8.465 2.400 11.170 2.560 ;
        RECT  10.820 1.960 10.980 2.220 ;
        RECT  10.815 0.620 10.975 1.745 ;
        RECT  8.805 2.060 10.820 2.220 ;
        RECT  10.540 0.620 10.815 0.780 ;
        RECT  10.695 1.280 10.815 1.745 ;
        RECT  10.365 1.585 10.695 1.745 ;
        RECT  10.280 0.560 10.540 0.780 ;
        RECT  9.795 1.170 10.475 1.330 ;
        RECT  10.095 1.585 10.365 1.850 ;
        RECT  9.520 1.690 10.095 1.850 ;
        RECT  9.795 0.570 10.025 0.730 ;
        RECT  9.635 0.570 9.795 1.510 ;
        RECT  9.290 1.350 9.635 1.510 ;
        RECT  9.130 1.350 9.290 1.830 ;
        RECT  8.985 1.570 9.130 1.830 ;
        RECT  8.850 0.540 9.025 0.700 ;
        RECT  8.805 0.540 8.850 1.355 ;
        RECT  8.690 0.540 8.805 2.220 ;
        RECT  8.645 1.145 8.690 2.220 ;
        RECT  8.280 2.270 8.465 2.560 ;
        RECT  7.695 2.270 8.280 2.430 ;
        RECT  8.035 1.570 8.075 1.830 ;
        RECT  7.875 0.610 8.035 1.830 ;
        RECT  7.535 0.660 7.695 2.430 ;
        RECT  7.240 0.660 7.535 0.820 ;
        RECT  7.405 1.570 7.535 1.830 ;
        RECT  6.215 2.270 7.535 2.430 ;
        RECT  7.195 1.130 7.335 1.390 ;
        RECT  7.035 1.010 7.195 2.065 ;
        RECT  6.940 1.010 7.035 1.170 ;
        RECT  6.845 1.905 7.035 2.065 ;
        RECT  6.780 0.615 6.940 1.170 ;
        RECT  6.585 1.350 6.855 1.610 ;
        RECT  6.425 0.690 6.585 1.770 ;
        RECT  5.730 0.690 6.425 0.850 ;
        RECT  6.155 1.610 6.425 1.770 ;
        RECT  6.055 1.950 6.215 2.430 ;
        RECT  3.635 1.950 6.055 2.110 ;
        RECT  4.195 2.290 5.320 2.450 ;
        RECT  4.455 1.610 5.115 1.770 ;
        RECT  4.455 0.665 4.620 0.825 ;
        RECT  4.295 0.665 4.455 1.770 ;
        RECT  4.170 1.095 4.295 1.355 ;
        RECT  4.035 2.290 4.195 2.560 ;
        RECT  3.930 1.610 4.115 1.770 ;
        RECT  1.305 2.400 4.035 2.560 ;
        RECT  3.770 0.770 3.930 1.770 ;
        RECT  3.635 0.770 3.770 0.930 ;
        RECT  3.375 0.665 3.635 0.930 ;
        RECT  3.375 1.950 3.635 2.220 ;
        RECT  2.565 0.770 3.375 0.930 ;
        RECT  1.655 2.060 3.375 2.220 ;
        RECT  1.995 1.720 3.065 1.880 ;
        RECT  2.405 0.770 2.565 1.265 ;
        RECT  2.335 1.105 2.405 1.265 ;
        RECT  2.175 1.105 2.335 1.365 ;
        RECT  1.995 0.665 2.225 0.925 ;
        RECT  1.835 0.665 1.995 1.880 ;
        RECT  1.495 0.665 1.655 2.220 ;
        RECT  1.145 2.170 1.305 2.560 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.255 0.580 0.390 0.840 ;
        RECT  0.255 1.865 0.385 2.330 ;
        RECT  0.225 0.580 0.255 2.330 ;
        RECT  0.095 0.580 0.225 2.125 ;
    END
END SMDFFHQX1MTH

MACRO SMDFFHQX2MTH
    CLASS CORE ;
    FOREIGN SMDFFHQX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 17.630 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.205 1.185 1.465 ;
        RECT  0.920 1.205 1.130 1.990 ;
        END
        AntennaGateArea 0.0533 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 0.310 5.780 0.470 ;
        RECT  1.115 0.310 1.275 0.660 ;
        RECT  0.740 0.500 1.115 0.660 ;
        RECT  0.580 0.500 0.740 1.580 ;
        RECT  0.435 1.280 0.580 1.580 ;
        END
        AntennaGateArea 0.1469 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.985 1.230 6.245 1.420 ;
        RECT  5.640 1.260 5.985 1.420 ;
        RECT  5.430 1.260 5.640 1.580 ;
        RECT  4.810 1.260 5.430 1.420 ;
        RECT  4.650 1.160 4.810 1.420 ;
        END
        AntennaGateArea 0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.475 1.290 17.530 1.580 ;
        RECT  17.295 0.425 17.475 2.285 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 1.175 3.635 1.580 ;
        RECT  2.685 1.175 3.350 1.435 ;
        END
        AntennaGateArea 0.0884 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.375 0.470 8.510 0.770 ;
        RECT  8.215 0.470 8.375 1.250 ;
        END
        AntennaGateArea 0.0871 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.180 0.680 9.450 1.170 ;
        RECT  9.030 0.880 9.180 1.170 ;
        END
        AntennaGateArea 0.1417 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.945 -0.130 17.630 0.130 ;
        RECT  16.785 -0.130 16.945 1.025 ;
        RECT  15.975 -0.130 16.785 0.130 ;
        RECT  15.375 -0.130 15.975 0.300 ;
        RECT  13.580 -0.130 15.375 0.130 ;
        RECT  13.080 -0.130 13.580 0.300 ;
        RECT  11.215 -0.130 13.080 0.130 ;
        RECT  10.955 -0.130 11.215 0.300 ;
        RECT  10.545 -0.130 10.955 0.130 ;
        RECT  10.285 -0.130 10.545 0.300 ;
        RECT  9.465 -0.130 10.285 0.130 ;
        RECT  9.205 -0.130 9.465 0.300 ;
        RECT  7.190 -0.130 9.205 0.130 ;
        RECT  6.350 -0.130 7.190 0.300 ;
        RECT  0.840 -0.130 6.350 0.130 ;
        RECT  0.340 -0.130 0.840 0.300 ;
        RECT  0.000 -0.130 0.340 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.945 2.740 17.630 3.000 ;
        RECT  16.785 1.775 16.945 3.000 ;
        RECT  16.315 2.740 16.785 3.000 ;
        RECT  15.715 2.450 16.315 3.000 ;
        RECT  8.050 2.740 15.715 3.000 ;
        RECT  7.450 2.620 8.050 3.000 ;
        RECT  6.375 2.740 7.450 3.000 ;
        RECT  5.435 2.620 6.375 3.000 ;
        RECT  4.695 2.740 5.435 3.000 ;
        RECT  4.435 2.620 4.695 3.000 ;
        RECT  0.755 2.740 4.435 3.000 ;
        RECT  0.255 2.570 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.380 0.565 16.540 2.145 ;
        RECT  16.225 0.565 16.380 0.725 ;
        RECT  16.275 1.725 16.380 2.145 ;
        RECT  15.765 1.725 16.275 1.885 ;
        RECT  16.030 1.010 16.190 1.290 ;
        RECT  15.305 1.130 16.030 1.290 ;
        RECT  15.505 1.560 15.765 1.885 ;
        RECT  15.145 0.595 15.305 1.875 ;
        RECT  15.185 2.365 15.285 2.525 ;
        RECT  15.025 2.060 15.185 2.525 ;
        RECT  14.860 0.595 15.145 0.755 ;
        RECT  14.600 1.715 15.145 1.875 ;
        RECT  14.415 2.060 15.025 2.220 ;
        RECT  14.685 0.935 14.945 1.195 ;
        RECT  14.600 0.495 14.860 0.755 ;
        RECT  11.675 2.400 14.805 2.560 ;
        RECT  14.415 1.035 14.685 1.195 ;
        RECT  14.255 1.035 14.415 2.220 ;
        RECT  12.015 2.060 14.255 2.220 ;
        RECT  14.070 0.580 14.170 0.840 ;
        RECT  13.910 0.580 14.070 1.875 ;
        RECT  13.250 0.680 13.910 0.840 ;
        RECT  13.775 1.715 13.910 1.875 ;
        RECT  13.595 1.120 13.730 1.380 ;
        RECT  13.435 1.120 13.595 1.610 ;
        RECT  12.910 1.450 13.435 1.610 ;
        RECT  13.090 0.680 13.250 1.265 ;
        RECT  12.750 0.650 12.910 1.610 ;
        RECT  12.355 0.650 12.750 0.810 ;
        RECT  12.355 1.450 12.750 1.610 ;
        RECT  12.015 1.010 12.555 1.270 ;
        RECT  12.195 0.550 12.355 0.810 ;
        RECT  12.195 1.450 12.355 1.880 ;
        RECT  11.855 0.635 12.015 2.220 ;
        RECT  10.975 0.635 11.855 0.795 ;
        RECT  11.515 1.000 11.675 2.560 ;
        RECT  11.365 1.000 11.515 1.160 ;
        RECT  10.980 1.960 11.515 2.120 ;
        RECT  11.175 2.300 11.335 2.560 ;
        RECT  8.465 2.400 11.175 2.560 ;
        RECT  10.975 1.310 11.075 1.470 ;
        RECT  10.820 1.960 10.980 2.220 ;
        RECT  10.815 0.635 10.975 1.745 ;
        RECT  8.805 2.060 10.820 2.220 ;
        RECT  10.545 0.635 10.815 0.795 ;
        RECT  10.365 1.585 10.815 1.745 ;
        RECT  10.285 0.585 10.545 0.795 ;
        RECT  9.795 1.170 10.475 1.330 ;
        RECT  10.095 1.585 10.365 1.850 ;
        RECT  9.520 1.690 10.095 1.850 ;
        RECT  9.795 0.540 10.035 0.700 ;
        RECT  9.635 0.540 9.795 1.510 ;
        RECT  9.290 1.350 9.635 1.510 ;
        RECT  9.130 1.350 9.290 1.795 ;
        RECT  8.985 1.535 9.130 1.795 ;
        RECT  8.850 0.540 8.995 0.700 ;
        RECT  8.805 0.540 8.850 1.355 ;
        RECT  8.690 0.540 8.805 2.220 ;
        RECT  8.645 1.145 8.690 2.220 ;
        RECT  8.280 2.270 8.465 2.560 ;
        RECT  7.695 2.270 8.280 2.430 ;
        RECT  8.035 1.570 8.075 1.830 ;
        RECT  7.875 0.610 8.035 1.830 ;
        RECT  7.535 0.660 7.695 2.430 ;
        RECT  7.240 0.660 7.535 0.820 ;
        RECT  7.405 1.570 7.535 1.830 ;
        RECT  5.680 2.270 7.535 2.430 ;
        RECT  7.195 1.130 7.335 1.390 ;
        RECT  7.035 1.010 7.195 2.065 ;
        RECT  6.940 1.010 7.035 1.170 ;
        RECT  6.845 1.905 7.035 2.065 ;
        RECT  6.780 0.610 6.940 1.170 ;
        RECT  6.585 1.350 6.855 1.610 ;
        RECT  6.425 0.680 6.585 1.760 ;
        RECT  5.730 0.680 6.425 0.840 ;
        RECT  6.155 1.600 6.425 1.760 ;
        RECT  5.520 1.940 5.680 2.430 ;
        RECT  3.600 1.940 5.520 2.100 ;
        RECT  4.195 2.280 5.320 2.440 ;
        RECT  4.455 1.600 5.115 1.760 ;
        RECT  4.455 0.660 4.620 0.820 ;
        RECT  4.295 0.660 4.455 1.760 ;
        RECT  4.170 1.095 4.295 1.355 ;
        RECT  4.035 2.280 4.195 2.560 ;
        RECT  3.975 1.600 4.115 1.760 ;
        RECT  1.305 2.400 4.035 2.560 ;
        RECT  3.815 0.770 3.975 1.760 ;
        RECT  3.700 0.770 3.815 0.930 ;
        RECT  3.390 0.655 3.700 0.930 ;
        RECT  3.315 1.940 3.600 2.220 ;
        RECT  2.505 0.770 3.390 0.930 ;
        RECT  1.655 2.060 3.315 2.220 ;
        RECT  1.995 1.720 3.065 1.880 ;
        RECT  2.345 0.770 2.505 1.265 ;
        RECT  2.335 1.105 2.345 1.265 ;
        RECT  2.175 1.105 2.335 1.365 ;
        RECT  1.995 0.665 2.165 0.925 ;
        RECT  1.835 0.665 1.995 1.880 ;
        RECT  1.495 0.665 1.655 2.220 ;
        RECT  1.145 2.170 1.305 2.560 ;
        RECT  0.385 2.170 1.145 2.330 ;
        RECT  0.255 0.600 0.400 0.860 ;
        RECT  0.255 1.865 0.385 2.330 ;
        RECT  0.225 0.600 0.255 2.330 ;
        RECT  0.095 0.600 0.225 2.125 ;
    END
END SMDFFHQX2MTH

MACRO SMDFFHQX4MTH
    CLASS CORE ;
    FOREIGN SMDFFHQX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.040 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 1.270 1.185 1.990 ;
        RECT  0.920 1.700 0.950 1.990 ;
        END
        AntennaGateArea 0.0806 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 0.310 5.780 0.470 ;
        RECT  1.115 0.310 1.275 0.660 ;
        RECT  0.745 0.500 1.115 0.660 ;
        RECT  0.585 0.500 0.745 1.580 ;
        RECT  0.435 1.280 0.585 1.580 ;
        END
        AntennaGateArea 0.1599 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.985 1.230 6.245 1.420 ;
        RECT  5.640 1.260 5.985 1.420 ;
        RECT  5.430 1.260 5.640 1.580 ;
        RECT  4.810 1.260 5.430 1.420 ;
        RECT  4.650 1.160 4.810 1.420 ;
        END
        AntennaGateArea 0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  17.475 1.290 17.530 1.580 ;
        RECT  17.295 0.425 17.475 2.285 ;
        RECT  17.195 0.425 17.295 1.025 ;
        RECT  17.195 1.685 17.295 2.285 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 1.175 3.635 1.580 ;
        RECT  2.795 1.175 3.350 1.435 ;
        END
        AntennaGateArea 0.1599 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.375 0.470 8.510 0.760 ;
        RECT  8.215 0.470 8.375 1.250 ;
        END
        AntennaGateArea 0.1352 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.180 0.595 9.450 1.130 ;
        RECT  9.030 0.880 9.180 1.130 ;
        END
        AntennaGateArea 0.2015 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.865 -0.130 18.040 0.130 ;
        RECT  17.705 -0.130 17.865 1.025 ;
        RECT  16.840 -0.130 17.705 0.130 ;
        RECT  16.680 -0.130 16.840 1.025 ;
        RECT  16.305 -0.130 16.680 0.300 ;
        RECT  15.700 -0.130 16.305 0.130 ;
        RECT  15.480 -0.130 15.700 0.855 ;
        RECT  15.005 -0.130 15.480 0.300 ;
        RECT  13.615 -0.130 15.005 0.130 ;
        RECT  13.015 -0.130 13.615 0.300 ;
        RECT  11.315 -0.130 13.015 0.130 ;
        RECT  10.715 -0.130 11.315 0.300 ;
        RECT  6.850 -0.130 10.715 0.130 ;
        RECT  6.010 -0.130 6.850 0.300 ;
        RECT  0.765 -0.130 6.010 0.130 ;
        RECT  0.265 -0.130 0.765 0.300 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.865 2.740 18.040 3.000 ;
        RECT  17.705 1.775 17.865 3.000 ;
        RECT  16.825 2.740 17.705 3.000 ;
        RECT  16.305 2.450 16.825 3.000 ;
        RECT  16.115 2.740 16.305 3.000 ;
        RECT  15.595 2.450 16.115 3.000 ;
        RECT  8.050 2.740 15.595 3.000 ;
        RECT  7.450 2.620 8.050 3.000 ;
        RECT  6.375 2.740 7.450 3.000 ;
        RECT  5.435 2.620 6.375 3.000 ;
        RECT  4.790 2.740 5.435 3.000 ;
        RECT  4.530 2.620 4.790 3.000 ;
        RECT  0.755 2.740 4.530 3.000 ;
        RECT  0.255 2.570 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.315 0.645 16.475 2.145 ;
        RECT  16.115 0.645 16.315 0.805 ;
        RECT  16.205 1.725 16.315 2.145 ;
        RECT  15.575 1.725 16.205 1.885 ;
        RECT  15.965 1.190 16.125 1.450 ;
        RECT  15.180 1.190 15.965 1.350 ;
        RECT  15.415 1.560 15.575 1.885 ;
        RECT  15.205 2.365 15.305 2.525 ;
        RECT  15.045 2.060 15.205 2.525 ;
        RECT  15.020 0.565 15.180 1.875 ;
        RECT  14.435 2.060 15.045 2.220 ;
        RECT  14.745 0.565 15.020 0.725 ;
        RECT  14.615 1.715 15.020 1.875 ;
        RECT  11.855 2.400 14.825 2.560 ;
        RECT  14.485 0.465 14.745 0.725 ;
        RECT  14.435 1.035 14.535 1.195 ;
        RECT  14.275 1.035 14.435 2.220 ;
        RECT  12.195 2.060 14.275 2.220 ;
        RECT  14.090 0.580 14.235 0.840 ;
        RECT  13.975 0.580 14.090 1.875 ;
        RECT  13.930 0.680 13.975 1.875 ;
        RECT  13.270 0.680 13.930 0.840 ;
        RECT  13.795 1.715 13.930 1.875 ;
        RECT  13.610 1.190 13.750 1.450 ;
        RECT  13.450 1.190 13.610 1.765 ;
        RECT  12.930 1.605 13.450 1.765 ;
        RECT  13.110 0.680 13.270 1.265 ;
        RECT  12.770 0.655 12.930 1.765 ;
        RECT  12.590 0.655 12.770 0.815 ;
        RECT  12.620 1.605 12.770 1.765 ;
        RECT  12.460 1.605 12.620 1.865 ;
        RECT  12.430 0.555 12.590 0.815 ;
        RECT  12.195 1.005 12.590 1.265 ;
        RECT  12.035 0.620 12.195 2.220 ;
        RECT  11.035 0.620 12.035 0.780 ;
        RECT  11.695 1.035 11.855 2.560 ;
        RECT  11.375 1.035 11.695 1.195 ;
        RECT  10.980 1.960 11.695 2.120 ;
        RECT  8.465 2.400 11.515 2.560 ;
        RECT  10.875 0.620 11.035 1.745 ;
        RECT  10.820 1.960 10.980 2.220 ;
        RECT  10.435 0.620 10.875 0.780 ;
        RECT  10.305 1.585 10.875 1.745 ;
        RECT  8.850 2.060 10.820 2.220 ;
        RECT  9.795 1.170 10.475 1.330 ;
        RECT  10.175 0.520 10.435 0.780 ;
        RECT  10.045 1.585 10.305 1.880 ;
        RECT  9.675 1.720 10.045 1.880 ;
        RECT  9.795 0.465 9.925 0.625 ;
        RECT  9.635 0.465 9.795 1.495 ;
        RECT  9.245 1.335 9.635 1.495 ;
        RECT  9.045 1.335 9.245 1.595 ;
        RECT  8.850 0.415 8.945 0.675 ;
        RECT  8.690 0.415 8.850 2.220 ;
        RECT  8.280 2.270 8.465 2.560 ;
        RECT  7.695 2.270 8.280 2.430 ;
        RECT  8.035 1.645 8.075 1.905 ;
        RECT  7.875 0.415 8.035 1.905 ;
        RECT  7.535 0.615 7.695 2.430 ;
        RECT  7.240 0.615 7.535 0.775 ;
        RECT  7.405 1.660 7.535 1.920 ;
        RECT  6.215 2.270 7.535 2.430 ;
        RECT  7.195 1.185 7.335 1.445 ;
        RECT  7.035 1.010 7.195 2.065 ;
        RECT  6.940 1.010 7.035 1.170 ;
        RECT  6.845 1.905 7.035 2.065 ;
        RECT  6.780 0.615 6.940 1.170 ;
        RECT  6.585 1.350 6.855 1.610 ;
        RECT  6.425 0.760 6.585 1.760 ;
        RECT  5.990 0.760 6.425 0.920 ;
        RECT  6.155 1.600 6.425 1.760 ;
        RECT  6.055 1.940 6.215 2.430 ;
        RECT  3.605 1.940 6.055 2.100 ;
        RECT  5.730 0.680 5.990 0.920 ;
        RECT  3.950 2.280 5.320 2.440 ;
        RECT  4.455 1.600 5.115 1.760 ;
        RECT  4.455 0.665 4.660 0.825 ;
        RECT  4.295 0.665 4.455 1.760 ;
        RECT  4.210 1.095 4.295 1.360 ;
        RECT  4.170 1.095 4.210 1.355 ;
        RECT  3.975 0.665 4.115 0.915 ;
        RECT  3.975 1.600 4.115 1.760 ;
        RECT  3.855 0.665 3.975 1.760 ;
        RECT  3.790 2.280 3.950 2.560 ;
        RECT  3.815 0.770 3.855 1.760 ;
        RECT  2.615 0.770 3.815 0.930 ;
        RECT  1.245 2.400 3.790 2.560 ;
        RECT  3.345 1.940 3.605 2.220 ;
        RECT  1.655 2.060 3.345 2.220 ;
        RECT  1.995 1.720 3.065 1.880 ;
        RECT  2.455 0.770 2.615 1.265 ;
        RECT  2.335 1.105 2.455 1.265 ;
        RECT  2.175 1.105 2.335 1.365 ;
        RECT  1.995 0.650 2.275 0.860 ;
        RECT  1.835 0.650 1.995 1.880 ;
        RECT  1.495 0.665 1.655 2.220 ;
        RECT  1.085 2.170 1.245 2.560 ;
        RECT  0.385 2.170 1.085 2.330 ;
        RECT  0.255 0.555 0.405 0.870 ;
        RECT  0.255 1.865 0.385 2.330 ;
        RECT  0.225 0.555 0.255 2.330 ;
        RECT  0.095 0.555 0.225 2.125 ;
    END
END SMDFFHQX4MTH

MACRO SMDFFHQX8MTH
    CLASS CORE ;
    FOREIGN SMDFFHQX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 18.860 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SI
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.950 1.270 1.185 1.990 ;
        RECT  0.920 1.700 0.950 1.990 ;
        END
        AntennaGateArea 0.0806 ;
    END SI
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.275 0.310 5.780 0.470 ;
        RECT  1.115 0.310 1.275 0.660 ;
        RECT  0.745 0.500 1.115 0.660 ;
        RECT  0.585 0.500 0.745 1.580 ;
        RECT  0.435 1.280 0.585 1.580 ;
        END
        AntennaGateArea 0.1599 ;
    END SE
    PIN S0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.985 1.230 6.245 1.420 ;
        RECT  5.640 1.260 5.985 1.420 ;
        RECT  5.430 1.260 5.640 1.580 ;
        RECT  4.810 1.260 5.430 1.420 ;
        RECT  4.650 1.160 4.810 1.420 ;
        END
        AntennaGateArea 0.1235 ;
    END S0
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.265 1.685 18.335 2.285 ;
        RECT  18.005 0.425 18.265 2.285 ;
        RECT  17.265 1.290 18.005 1.580 ;
        RECT  17.245 1.290 17.265 2.285 ;
        RECT  16.985 0.425 17.245 2.285 ;
        END
        AntennaDiffArea 1.2 ;
    END Q
    PIN D1
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.350 1.175 3.635 1.580 ;
        RECT  2.795 1.175 3.350 1.435 ;
        END
        AntennaGateArea 0.1599 ;
    END D1
    PIN D0
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.375 0.470 8.510 0.760 ;
        RECT  8.215 0.470 8.375 1.250 ;
        END
        AntennaGateArea 0.1352 ;
    END D0
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.180 0.595 9.450 1.130 ;
        RECT  9.030 0.880 9.180 1.130 ;
        END
        AntennaGateArea 0.2015 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  18.685 -0.130 18.860 0.130 ;
        RECT  18.485 -0.130 18.685 1.025 ;
        RECT  17.685 -0.130 18.485 0.130 ;
        RECT  17.465 -0.130 17.685 1.025 ;
        RECT  16.605 -0.130 17.465 0.130 ;
        RECT  16.105 -0.130 16.605 0.300 ;
        RECT  15.660 -0.130 16.105 0.130 ;
        RECT  15.440 -0.130 15.660 0.855 ;
        RECT  15.005 -0.130 15.440 0.300 ;
        RECT  13.615 -0.130 15.005 0.130 ;
        RECT  13.015 -0.130 13.615 0.300 ;
        RECT  11.315 -0.130 13.015 0.130 ;
        RECT  10.715 -0.130 11.315 0.300 ;
        RECT  6.850 -0.130 10.715 0.130 ;
        RECT  6.010 -0.130 6.850 0.300 ;
        RECT  0.765 -0.130 6.010 0.130 ;
        RECT  0.265 -0.130 0.765 0.300 ;
        RECT  0.000 -0.130 0.265 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  17.805 2.740 18.860 3.000 ;
        RECT  17.585 1.770 17.805 3.000 ;
        RECT  16.775 2.740 17.585 3.000 ;
        RECT  16.170 2.450 16.775 3.000 ;
        RECT  15.985 2.740 16.170 3.000 ;
        RECT  15.720 2.450 15.985 3.000 ;
        RECT  8.050 2.740 15.720 3.000 ;
        RECT  7.450 2.620 8.050 3.000 ;
        RECT  6.375 2.740 7.450 3.000 ;
        RECT  5.435 2.620 6.375 3.000 ;
        RECT  4.685 2.740 5.435 3.000 ;
        RECT  4.425 2.620 4.685 3.000 ;
        RECT  0.755 2.740 4.425 3.000 ;
        RECT  0.255 2.570 0.755 3.000 ;
        RECT  0.000 2.740 0.255 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  16.305 0.645 16.465 2.145 ;
        RECT  16.020 0.645 16.305 0.805 ;
        RECT  16.195 1.725 16.305 2.145 ;
        RECT  15.565 1.725 16.195 1.885 ;
        RECT  15.930 1.190 16.090 1.450 ;
        RECT  15.180 1.190 15.930 1.350 ;
        RECT  15.405 1.560 15.565 1.885 ;
        RECT  15.205 2.365 15.305 2.525 ;
        RECT  15.045 2.060 15.205 2.525 ;
        RECT  15.020 0.565 15.180 1.875 ;
        RECT  14.435 2.060 15.045 2.220 ;
        RECT  14.745 0.565 15.020 0.725 ;
        RECT  14.615 1.715 15.020 1.875 ;
        RECT  11.855 2.400 14.825 2.560 ;
        RECT  14.485 0.465 14.745 0.725 ;
        RECT  14.435 1.035 14.535 1.195 ;
        RECT  14.275 1.035 14.435 2.220 ;
        RECT  12.195 2.060 14.275 2.220 ;
        RECT  14.090 0.580 14.235 0.840 ;
        RECT  13.975 0.580 14.090 1.875 ;
        RECT  13.930 0.680 13.975 1.875 ;
        RECT  13.270 0.680 13.930 0.840 ;
        RECT  13.795 1.715 13.930 1.875 ;
        RECT  13.610 1.190 13.750 1.450 ;
        RECT  13.450 1.190 13.610 1.765 ;
        RECT  12.930 1.605 13.450 1.765 ;
        RECT  13.110 0.680 13.270 1.265 ;
        RECT  12.770 0.655 12.930 1.765 ;
        RECT  12.590 0.655 12.770 0.815 ;
        RECT  12.620 1.605 12.770 1.765 ;
        RECT  12.460 1.605 12.620 1.865 ;
        RECT  12.430 0.555 12.590 0.815 ;
        RECT  12.195 1.005 12.590 1.265 ;
        RECT  12.035 0.620 12.195 2.220 ;
        RECT  11.035 0.620 12.035 0.780 ;
        RECT  11.695 1.035 11.855 2.560 ;
        RECT  11.375 1.035 11.695 1.195 ;
        RECT  10.980 1.960 11.695 2.120 ;
        RECT  8.465 2.400 11.515 2.560 ;
        RECT  10.875 0.620 11.035 1.745 ;
        RECT  10.820 1.960 10.980 2.220 ;
        RECT  10.435 0.620 10.875 0.780 ;
        RECT  10.305 1.585 10.875 1.745 ;
        RECT  8.850 2.060 10.820 2.220 ;
        RECT  9.795 1.170 10.475 1.330 ;
        RECT  10.175 0.520 10.435 0.780 ;
        RECT  10.045 1.585 10.305 1.880 ;
        RECT  9.675 1.720 10.045 1.880 ;
        RECT  9.795 0.465 9.925 0.625 ;
        RECT  9.635 0.465 9.795 1.495 ;
        RECT  9.245 1.335 9.635 1.495 ;
        RECT  9.045 1.335 9.245 1.595 ;
        RECT  8.850 0.415 8.945 0.675 ;
        RECT  8.690 0.415 8.850 2.220 ;
        RECT  8.280 2.270 8.465 2.560 ;
        RECT  7.695 2.270 8.280 2.430 ;
        RECT  8.035 1.645 8.075 1.905 ;
        RECT  7.875 0.415 8.035 1.905 ;
        RECT  7.535 0.615 7.695 2.430 ;
        RECT  7.240 0.615 7.535 0.775 ;
        RECT  7.405 1.660 7.535 1.920 ;
        RECT  6.215 2.270 7.535 2.430 ;
        RECT  7.195 1.185 7.335 1.445 ;
        RECT  7.035 1.010 7.195 2.065 ;
        RECT  6.940 1.010 7.035 1.170 ;
        RECT  6.845 1.905 7.035 2.065 ;
        RECT  6.780 0.615 6.940 1.170 ;
        RECT  6.585 1.350 6.855 1.610 ;
        RECT  6.425 0.760 6.585 1.760 ;
        RECT  5.990 0.760 6.425 0.920 ;
        RECT  6.155 1.600 6.425 1.760 ;
        RECT  6.055 1.940 6.215 2.430 ;
        RECT  3.605 1.940 6.055 2.100 ;
        RECT  5.730 0.680 5.990 0.920 ;
        RECT  3.950 2.280 5.320 2.440 ;
        RECT  4.455 1.600 5.115 1.760 ;
        RECT  4.455 0.665 4.660 0.825 ;
        RECT  4.295 0.665 4.455 1.760 ;
        RECT  4.210 1.095 4.295 1.360 ;
        RECT  4.170 1.095 4.210 1.355 ;
        RECT  3.975 0.665 4.115 0.915 ;
        RECT  3.975 1.600 4.115 1.760 ;
        RECT  3.855 0.665 3.975 1.760 ;
        RECT  3.790 2.280 3.950 2.560 ;
        RECT  3.815 0.770 3.855 1.760 ;
        RECT  2.615 0.770 3.815 0.930 ;
        RECT  1.245 2.400 3.790 2.560 ;
        RECT  3.345 1.940 3.605 2.220 ;
        RECT  1.655 2.060 3.345 2.220 ;
        RECT  1.995 1.720 3.065 1.880 ;
        RECT  2.455 0.770 2.615 1.265 ;
        RECT  2.335 1.105 2.455 1.265 ;
        RECT  2.175 1.105 2.335 1.365 ;
        RECT  1.995 0.650 2.275 0.860 ;
        RECT  1.835 0.650 1.995 1.880 ;
        RECT  1.495 0.665 1.655 2.220 ;
        RECT  1.085 2.170 1.245 2.560 ;
        RECT  0.385 2.170 1.085 2.330 ;
        RECT  0.255 0.555 0.405 0.870 ;
        RECT  0.255 1.865 0.385 2.330 ;
        RECT  0.225 0.555 0.255 2.330 ;
        RECT  0.095 0.555 0.225 2.125 ;
    END
END SMDFFHQX8MTH

MACRO TBUFX12MTH
    CLASS CORE ;
    FOREIGN TBUFX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  6.075 0.390 6.335 2.285 ;
        RECT  5.315 0.975 6.075 1.745 ;
        RECT  5.055 0.360 5.315 2.450 ;
        RECT  4.785 0.745 5.055 2.125 ;
        RECT  4.305 0.745 4.785 1.255 ;
        RECT  4.285 1.805 4.785 2.125 ;
        RECT  4.295 0.745 4.305 0.945 ;
        RECT  4.035 0.410 4.295 0.945 ;
        RECT  4.025 1.805 4.285 2.450 ;
        END
        AntennaDiffArea 1.731 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.080 0.505 1.680 ;
        END
        AntennaGateArea 0.2938 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.170 3.260 1.430 ;
        RECT  2.560 1.170 2.770 1.580 ;
        END
        AntennaGateArea 0.5265 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 -0.130 6.970 0.130 ;
        RECT  6.585 -0.130 6.845 0.985 ;
        RECT  5.825 -0.130 6.585 0.130 ;
        RECT  5.565 -0.130 5.825 0.795 ;
        RECT  4.805 -0.130 5.565 0.130 ;
        RECT  4.545 -0.130 4.805 0.565 ;
        RECT  0.815 -0.130 4.545 0.130 ;
        RECT  0.215 -0.130 0.815 0.300 ;
        RECT  0.000 -0.130 0.215 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 2.740 6.970 3.000 ;
        RECT  6.585 1.800 6.845 3.000 ;
        RECT  5.825 2.740 6.585 3.000 ;
        RECT  5.565 1.925 5.825 3.000 ;
        RECT  4.795 2.740 5.565 3.000 ;
        RECT  4.535 2.305 4.795 3.000 ;
        RECT  0.545 2.740 4.535 3.000 ;
        RECT  0.285 2.570 0.545 3.000 ;
        RECT  0.000 2.740 0.285 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.345 1.435 4.605 1.625 ;
        RECT  3.845 1.465 4.345 1.625 ;
        RECT  3.755 1.125 4.125 1.285 ;
        RECT  3.685 1.465 3.845 1.920 ;
        RECT  3.595 0.765 3.755 1.285 ;
        RECT  3.345 1.760 3.685 1.920 ;
        RECT  3.345 0.765 3.595 0.925 ;
        RECT  3.085 0.665 3.345 0.925 ;
        RECT  3.085 1.760 3.345 2.360 ;
        RECT  2.375 0.765 3.085 0.925 ;
        RECT  2.415 1.760 3.085 1.920 ;
        RECT  2.315 1.760 2.415 2.360 ;
        RECT  2.275 0.665 2.375 0.925 ;
        RECT  2.155 1.305 2.315 2.360 ;
        RECT  2.115 0.310 2.275 0.925 ;
        RECT  1.865 1.305 2.155 1.465 ;
        RECT  1.355 2.060 2.155 2.220 ;
        RECT  1.425 0.310 2.115 0.470 ;
        RECT  1.645 1.645 1.905 1.880 ;
        RECT  1.705 0.670 1.865 1.465 ;
        RECT  1.605 0.670 1.705 0.930 ;
        RECT  1.425 1.645 1.645 1.805 ;
        RECT  0.885 2.400 1.615 2.560 ;
        RECT  1.265 0.310 1.425 1.805 ;
        RECT  1.095 2.030 1.355 2.220 ;
        RECT  1.095 0.590 1.265 0.830 ;
        RECT  0.885 1.010 1.085 1.270 ;
        RECT  0.725 0.615 0.885 2.560 ;
        RECT  0.120 0.615 0.725 0.855 ;
        RECT  0.165 1.980 0.725 2.240 ;
    END
END TBUFX12MTH

MACRO TBUFX16MTH
    CLASS CORE ;
    FOREIGN TBUFX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.790 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  6.945 0.345 7.645 2.465 ;
        RECT  6.245 0.885 6.945 1.965 ;
        RECT  5.040 0.350 6.245 2.520 ;
        RECT  4.125 0.350 5.040 0.945 ;
        RECT  4.110 1.865 5.040 2.520 ;
        END
        AntennaDiffArea 2.331 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.355 1.515 ;
        END
        AntennaGateArea 0.3822 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.135 3.060 1.580 ;
        END
        AntennaGateArea 0.611 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.755 -0.130 7.790 0.130 ;
        RECT  6.495 -0.130 6.755 0.705 ;
        RECT  3.875 -0.130 6.495 0.130 ;
        RECT  3.615 -0.130 3.875 0.945 ;
        RECT  2.855 -0.130 3.615 0.130 ;
        RECT  2.595 -0.130 2.855 0.605 ;
        RECT  0.000 -0.130 2.595 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.755 2.740 7.790 3.000 ;
        RECT  6.495 2.145 6.755 3.000 ;
        RECT  0.720 2.740 6.495 3.000 ;
        RECT  0.125 2.570 0.720 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.450 1.385 4.710 1.685 ;
        RECT  3.430 1.525 4.450 1.685 ;
        RECT  3.430 1.125 4.215 1.285 ;
        RECT  3.365 0.785 3.430 1.285 ;
        RECT  3.270 1.525 3.430 2.360 ;
        RECT  3.270 0.435 3.365 1.285 ;
        RECT  3.105 0.435 3.270 0.945 ;
        RECT  3.170 1.760 3.270 2.360 ;
        RECT  2.500 1.760 3.170 1.920 ;
        RECT  2.335 0.785 3.105 0.945 ;
        RECT  2.365 1.760 2.500 2.260 ;
        RECT  2.240 1.255 2.365 2.260 ;
        RECT  2.095 0.310 2.335 0.945 ;
        RECT  2.205 1.255 2.240 2.220 ;
        RECT  1.785 1.255 2.205 1.415 ;
        RECT  1.400 2.060 2.205 2.220 ;
        RECT  1.445 0.310 2.095 0.470 ;
        RECT  1.730 1.595 1.990 1.880 ;
        RECT  1.625 0.655 1.785 1.415 ;
        RECT  1.445 1.595 1.730 1.755 ;
        RECT  1.060 2.400 1.710 2.560 ;
        RECT  1.285 0.310 1.445 1.755 ;
        RECT  1.240 1.935 1.400 2.220 ;
        RECT  1.065 0.545 1.285 0.805 ;
        RECT  0.900 1.075 1.060 2.560 ;
        RECT  0.885 1.075 0.900 1.335 ;
        RECT  0.125 1.860 0.900 2.120 ;
        RECT  0.725 0.410 0.885 1.335 ;
        RECT  0.125 0.410 0.725 0.570 ;
    END
END TBUFX16MTH

MACRO TBUFX1MTH
    CLASS CORE ;
    FOREIGN TBUFX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.430 0.475 3.590 2.310 ;
        RECT  3.190 0.475 3.430 0.735 ;
        RECT  3.380 1.700 3.430 2.310 ;
        RECT  3.195 2.050 3.380 2.310 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.195 0.510 1.460 ;
        RECT  0.100 1.195 0.310 1.580 ;
        END
        AntennaGateArea 0.1079 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.050 1.630 2.415 1.990 ;
        END
        AntennaGateArea 0.0546 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 -0.130 3.690 0.130 ;
        RECT  2.650 -0.130 2.910 0.740 ;
        RECT  1.010 -0.130 2.650 0.130 ;
        RECT  0.410 -0.130 1.010 0.485 ;
        RECT  0.000 -0.130 0.410 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 2.740 3.690 3.000 ;
        RECT  2.680 2.185 2.940 3.000 ;
        RECT  0.385 2.740 2.680 3.000 ;
        RECT  0.145 2.250 0.385 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.090 0.920 3.250 1.315 ;
        RECT  2.440 0.920 3.090 1.080 ;
        RECT  2.595 1.290 2.855 1.695 ;
        RECT  2.100 1.290 2.595 1.450 ;
        RECT  2.280 0.405 2.440 1.080 ;
        RECT  1.870 2.215 2.360 2.555 ;
        RECT  1.570 0.405 2.280 0.595 ;
        RECT  1.940 0.885 2.100 1.450 ;
        RECT  1.870 1.290 1.940 1.450 ;
        RECT  1.710 1.290 1.870 2.555 ;
        RECT  0.975 2.395 1.710 2.555 ;
        RECT  1.530 0.405 1.570 1.025 ;
        RECT  1.370 0.405 1.530 2.210 ;
        RECT  1.325 1.950 1.370 2.210 ;
        RECT  1.000 0.700 1.160 0.975 ;
        RECT  0.875 1.805 1.145 2.080 ;
        RECT  0.875 0.815 1.000 0.975 ;
        RECT  0.715 2.305 0.975 2.555 ;
        RECT  0.715 0.815 0.875 2.080 ;
        RECT  0.125 0.815 0.715 0.975 ;
        RECT  0.605 1.685 0.715 2.080 ;
    END
END TBUFX1MTH

MACRO TBUFX20MTH
    CLASS CORE ;
    FOREIGN TBUFX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  9.695 0.355 10.095 2.355 ;
        RECT  9.075 0.840 9.695 1.785 ;
        RECT  8.055 0.350 9.075 2.520 ;
        RECT  5.915 0.350 8.055 0.905 ;
        RECT  5.885 1.845 8.055 2.520 ;
        END
        AntennaDiffArea 2.881 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.405 1.505 ;
        END
        AntennaGateArea 0.4628 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.000 1.225 4.535 1.485 ;
        RECT  3.695 1.225 4.000 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 -0.130 10.660 0.130 ;
        RECT  10.275 -0.130 10.535 0.995 ;
        RECT  9.515 -0.130 10.275 0.130 ;
        RECT  9.255 -0.130 9.515 0.660 ;
        RECT  5.635 -0.130 9.255 0.130 ;
        RECT  5.375 -0.130 5.635 0.495 ;
        RECT  3.795 -0.130 5.375 0.130 ;
        RECT  3.535 -0.130 3.795 0.640 ;
        RECT  1.865 -0.130 3.535 0.130 ;
        RECT  1.605 -0.130 1.865 0.300 ;
        RECT  0.000 -0.130 1.605 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.535 2.740 10.660 3.000 ;
        RECT  10.275 1.845 10.535 3.000 ;
        RECT  9.515 2.740 10.275 3.000 ;
        RECT  9.255 1.965 9.515 3.000 ;
        RECT  5.605 2.740 9.255 3.000 ;
        RECT  5.345 2.245 5.605 3.000 ;
        RECT  3.765 2.740 5.345 3.000 ;
        RECT  3.505 2.105 3.765 3.000 ;
        RECT  1.665 2.740 3.505 3.000 ;
        RECT  0.725 2.485 1.665 3.000 ;
        RECT  0.000 2.740 0.725 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.530 1.435 7.470 1.625 ;
        RECT  5.460 1.465 6.530 1.625 ;
        RECT  5.530 1.125 6.345 1.285 ;
        RECT  5.370 0.820 5.530 1.285 ;
        RECT  5.300 1.465 5.460 1.920 ;
        RECT  5.235 0.820 5.370 0.980 ;
        RECT  5.205 1.760 5.300 1.920 ;
        RECT  4.975 0.720 5.235 0.980 ;
        RECT  4.945 1.760 5.205 2.020 ;
        RECT  4.305 0.820 4.975 0.980 ;
        RECT  4.275 1.760 4.945 1.920 ;
        RECT  4.045 0.380 4.305 0.980 ;
        RECT  4.015 1.760 4.275 2.420 ;
        RECT  3.335 0.820 4.045 0.980 ;
        RECT  3.255 1.760 4.015 1.920 ;
        RECT  3.175 0.310 3.335 0.980 ;
        RECT  3.155 1.720 3.255 2.360 ;
        RECT  3.025 0.310 3.175 0.565 ;
        RECT  2.995 1.720 3.155 2.560 ;
        RECT  2.215 0.310 3.025 0.470 ;
        RECT  2.965 1.720 2.995 1.880 ;
        RECT  2.235 2.400 2.995 2.560 ;
        RECT  2.805 0.735 2.965 1.880 ;
        RECT  2.515 0.735 2.805 0.895 ;
        RECT  2.625 2.060 2.745 2.220 ;
        RECT  2.465 1.075 2.625 2.220 ;
        RECT  2.215 1.075 2.465 1.235 ;
        RECT  1.875 1.430 2.285 1.600 ;
        RECT  1.975 1.860 2.235 2.560 ;
        RECT  2.055 0.310 2.215 1.235 ;
        RECT  1.325 0.525 2.055 0.685 ;
        RECT  1.325 1.860 1.975 2.020 ;
        RECT  1.715 0.965 1.875 1.600 ;
        RECT  1.495 0.965 1.715 1.125 ;
        RECT  0.745 0.865 1.495 1.125 ;
        RECT  1.065 0.425 1.325 0.685 ;
        RECT  1.065 1.860 1.325 2.120 ;
        RECT  0.585 0.430 0.745 1.845 ;
        RECT  0.125 0.430 0.585 0.690 ;
        RECT  0.385 1.685 0.585 1.845 ;
        RECT  0.125 1.685 0.385 2.285 ;
    END
END TBUFX20MTH

MACRO TBUFX24MTH
    CLASS CORE ;
    FOREIGN TBUFX24MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 12.710 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  11.815 0.355 12.075 2.285 ;
        RECT  11.145 0.785 11.815 1.985 ;
        RECT  11.135 0.355 11.145 1.985 ;
        RECT  10.885 0.355 11.135 2.285 ;
        RECT  10.875 0.785 10.885 2.285 ;
        RECT  10.205 0.785 10.875 1.985 ;
        RECT  10.125 0.785 10.205 2.285 ;
        RECT  9.945 0.355 10.125 2.285 ;
        RECT  9.865 0.355 9.945 1.985 ;
        RECT  9.195 0.785 9.865 1.985 ;
        RECT  9.185 0.355 9.195 1.985 ;
        RECT  8.935 0.355 9.185 2.520 ;
        RECT  8.415 0.745 8.935 2.520 ;
        RECT  8.245 0.745 8.415 1.215 ;
        RECT  7.065 1.845 8.415 2.520 ;
        RECT  7.795 0.350 8.245 1.215 ;
        RECT  6.985 0.350 7.795 0.945 ;
        END
        AntennaDiffArea 3.481 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.355 1.665 ;
        END
        AntennaGateArea 0.5915 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.230 1.225 5.495 1.485 ;
        RECT  5.020 1.225 5.230 1.580 ;
        RECT  4.315 1.225 5.020 1.485 ;
        END
        AntennaGateArea 1.027 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.585 -0.130 12.710 0.130 ;
        RECT  12.325 -0.130 12.585 0.970 ;
        RECT  10.635 -0.130 12.325 0.130 ;
        RECT  10.375 -0.130 10.635 0.605 ;
        RECT  8.685 -0.130 10.375 0.130 ;
        RECT  8.425 -0.130 8.685 0.565 ;
        RECT  6.735 -0.130 8.425 0.130 ;
        RECT  6.475 -0.130 6.735 0.945 ;
        RECT  5.715 -0.130 6.475 0.130 ;
        RECT  5.455 -0.130 5.715 0.640 ;
        RECT  4.695 -0.130 5.455 0.130 ;
        RECT  4.435 -0.130 4.695 0.640 ;
        RECT  1.925 -0.130 4.435 0.130 ;
        RECT  1.765 -0.130 1.925 0.695 ;
        RECT  0.925 -0.130 1.765 0.130 ;
        RECT  0.665 -0.130 0.925 0.330 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.585 2.740 12.710 3.000 ;
        RECT  12.325 1.825 12.585 3.000 ;
        RECT  9.695 2.740 12.325 3.000 ;
        RECT  9.435 2.165 9.695 3.000 ;
        RECT  6.815 2.740 9.435 3.000 ;
        RECT  6.555 1.815 6.815 3.000 ;
        RECT  4.865 2.740 6.555 3.000 ;
        RECT  4.605 2.100 4.865 3.000 ;
        RECT  3.845 2.740 4.605 3.000 ;
        RECT  3.585 2.045 3.845 3.000 ;
        RECT  0.385 2.740 3.585 3.000 ;
        RECT  0.125 1.875 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.635 1.435 8.235 1.625 ;
        RECT  6.305 1.465 7.635 1.625 ;
        RECT  6.225 1.125 7.415 1.285 ;
        RECT  6.145 1.465 6.305 2.420 ;
        RECT  6.065 0.380 6.225 1.285 ;
        RECT  6.045 1.760 6.145 2.420 ;
        RECT  5.965 0.380 6.065 0.980 ;
        RECT  5.375 1.760 6.045 1.920 ;
        RECT  5.205 0.820 5.965 0.980 ;
        RECT  5.115 1.760 5.375 2.420 ;
        RECT  4.945 0.380 5.205 0.980 ;
        RECT  4.355 1.760 5.115 1.920 ;
        RECT  4.135 0.820 4.945 0.980 ;
        RECT  4.095 1.705 4.355 2.255 ;
        RECT  3.975 0.310 4.135 0.980 ;
        RECT  3.285 1.705 4.095 1.865 ;
        RECT  3.165 0.310 3.975 0.470 ;
        RECT  3.415 0.650 3.675 0.915 ;
        RECT  3.285 0.755 3.415 0.915 ;
        RECT  3.125 0.755 3.285 2.420 ;
        RECT  2.905 0.310 3.165 0.575 ;
        RECT  2.605 0.755 3.125 0.915 ;
        RECT  2.315 2.260 3.125 2.420 ;
        RECT  2.265 0.310 2.905 0.470 ;
        RECT  2.565 1.655 2.825 2.075 ;
        RECT  2.445 0.650 2.605 0.915 ;
        RECT  2.265 1.655 2.565 1.815 ;
        RECT  2.055 1.995 2.315 2.420 ;
        RECT  2.105 0.310 2.265 1.815 ;
        RECT  1.465 0.875 2.105 1.035 ;
        RECT  1.805 1.655 2.105 1.815 ;
        RECT  1.295 2.260 2.055 2.420 ;
        RECT  0.725 1.215 1.925 1.475 ;
        RECT  1.545 1.655 1.805 2.075 ;
        RECT  1.305 0.440 1.465 1.035 ;
        RECT  1.205 0.440 1.305 0.700 ;
        RECT  1.135 1.735 1.295 2.420 ;
        RECT  1.035 1.735 1.135 1.995 ;
        RECT  0.725 2.220 0.895 2.480 ;
        RECT  0.565 0.540 0.725 2.480 ;
        RECT  0.385 0.540 0.565 0.700 ;
        RECT  0.125 0.440 0.385 0.700 ;
    END
END TBUFX24MTH

MACRO TBUFX2MTH
    CLASS CORE ;
    FOREIGN TBUFX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.690 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.430 0.465 3.590 2.485 ;
        RECT  3.190 0.465 3.430 0.725 ;
        RECT  3.380 1.700 3.430 2.485 ;
        RECT  3.195 1.885 3.380 2.485 ;
        END
        AntennaDiffArea 0.449 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.195 0.510 1.460 ;
        RECT  0.100 1.195 0.310 1.580 ;
        END
        AntennaGateArea 0.1079 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.050 1.630 2.415 1.990 ;
        END
        AntennaGateArea 0.0871 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 -0.130 3.690 0.130 ;
        RECT  2.650 -0.130 2.910 0.765 ;
        RECT  1.010 -0.130 2.650 0.130 ;
        RECT  0.410 -0.130 1.010 0.485 ;
        RECT  0.000 -0.130 0.410 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.940 2.740 3.690 3.000 ;
        RECT  2.680 2.215 2.940 3.000 ;
        RECT  0.385 2.740 2.680 3.000 ;
        RECT  0.145 2.250 0.385 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.050 0.945 3.250 1.315 ;
        RECT  2.440 0.945 3.050 1.105 ;
        RECT  2.595 1.290 2.855 1.695 ;
        RECT  2.100 1.290 2.595 1.450 ;
        RECT  2.280 0.405 2.440 1.105 ;
        RECT  1.870 2.215 2.400 2.555 ;
        RECT  2.110 0.405 2.280 0.605 ;
        RECT  1.600 0.405 2.110 0.565 ;
        RECT  1.940 0.865 2.100 1.450 ;
        RECT  1.870 1.290 1.940 1.450 ;
        RECT  1.710 1.290 1.870 2.555 ;
        RECT  0.975 2.395 1.710 2.555 ;
        RECT  1.530 0.405 1.600 1.005 ;
        RECT  1.370 0.405 1.530 2.210 ;
        RECT  1.325 1.950 1.370 2.210 ;
        RECT  1.000 0.705 1.160 0.975 ;
        RECT  0.875 1.805 1.145 2.080 ;
        RECT  0.875 0.815 1.000 0.975 ;
        RECT  0.715 2.305 0.975 2.555 ;
        RECT  0.715 0.815 0.875 2.080 ;
        RECT  0.125 0.815 0.715 0.975 ;
        RECT  0.605 1.685 0.715 2.080 ;
    END
END TBUFX2MTH

MACRO TBUFX3MTH
    CLASS CORE ;
    FOREIGN TBUFX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.540 1.285 3.590 1.580 ;
        RECT  3.380 0.470 3.540 2.515 ;
        RECT  3.195 0.470 3.380 0.730 ;
        RECT  3.200 1.915 3.380 2.515 ;
        END
        AntennaDiffArea 0.452 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.195 0.535 1.460 ;
        RECT  0.100 1.195 0.310 1.580 ;
        END
        AntennaGateArea 0.1144 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.690 2.575 1.990 ;
        END
        AntennaGateArea 0.13 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.975 -0.130 4.100 0.130 ;
        RECT  3.720 -0.130 3.975 0.725 ;
        RECT  2.910 -0.130 3.720 0.130 ;
        RECT  2.650 -0.130 2.910 0.735 ;
        RECT  1.010 -0.130 2.650 0.130 ;
        RECT  0.410 -0.130 1.010 0.485 ;
        RECT  0.000 -0.130 0.410 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 2.740 4.100 3.000 ;
        RECT  3.760 1.915 3.970 3.000 ;
        RECT  2.940 2.740 3.760 3.000 ;
        RECT  2.680 2.210 2.940 3.000 ;
        RECT  0.385 2.740 2.680 3.000 ;
        RECT  0.145 2.250 0.385 3.000 ;
        RECT  0.000 2.740 0.145 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  2.940 0.920 3.200 1.170 ;
        RECT  2.940 1.350 3.200 1.730 ;
        RECT  2.470 0.920 2.940 1.080 ;
        RECT  2.100 1.350 2.940 1.510 ;
        RECT  2.310 0.425 2.470 1.080 ;
        RECT  1.925 2.170 2.400 2.430 ;
        RECT  1.570 0.425 2.310 0.615 ;
        RECT  1.940 1.025 2.100 1.510 ;
        RECT  1.925 1.350 1.940 1.510 ;
        RECT  1.765 1.350 1.925 2.550 ;
        RECT  0.955 2.390 1.765 2.550 ;
        RECT  1.530 0.425 1.570 1.025 ;
        RECT  1.370 0.425 1.530 2.210 ;
        RECT  1.325 1.950 1.370 2.210 ;
        RECT  1.000 0.705 1.160 0.975 ;
        RECT  0.875 1.805 1.145 2.085 ;
        RECT  0.875 0.815 1.000 0.975 ;
        RECT  0.695 2.305 0.955 2.550 ;
        RECT  0.715 0.815 0.875 2.085 ;
        RECT  0.125 0.815 0.715 0.975 ;
        RECT  0.605 1.685 0.715 2.085 ;
    END
END TBUFX3MTH

MACRO TBUFX4MTH
    CLASS CORE ;
    FOREIGN TBUFX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  3.790 0.910 4.000 2.025 ;
        RECT  3.465 0.910 3.790 1.090 ;
        RECT  3.460 1.845 3.790 2.025 ;
        RECT  3.285 0.475 3.465 1.090 ;
        RECT  3.200 1.845 3.460 2.450 ;
        RECT  3.195 0.475 3.285 0.735 ;
        END
        AntennaDiffArea 0.554 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.240 0.820 1.500 ;
        RECT  0.100 1.240 0.310 1.580 ;
        END
        AntennaGateArea 0.1235 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.280 2.570 1.580 ;
        END
        AntennaGateArea 0.1755 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.970 -0.130 4.100 0.130 ;
        RECT  3.715 -0.130 3.970 0.725 ;
        RECT  2.940 -0.130 3.715 0.130 ;
        RECT  2.680 -0.130 2.940 0.665 ;
        RECT  1.010 -0.130 2.680 0.130 ;
        RECT  0.410 -0.130 1.010 0.485 ;
        RECT  0.000 -0.130 0.410 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.980 2.740 4.100 3.000 ;
        RECT  3.715 2.215 3.980 3.000 ;
        RECT  2.935 2.740 3.715 3.000 ;
        RECT  2.670 2.210 2.935 3.000 ;
        RECT  0.385 2.740 2.670 3.000 ;
        RECT  0.135 2.250 0.385 3.000 ;
        RECT  0.000 2.740 0.135 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.285 1.395 3.545 1.655 ;
        RECT  2.920 1.495 3.285 1.655 ;
        RECT  2.800 0.940 3.060 1.295 ;
        RECT  2.760 1.495 2.920 1.920 ;
        RECT  2.400 0.940 2.800 1.100 ;
        RECT  2.400 1.760 2.760 1.920 ;
        RECT  2.240 0.405 2.400 1.100 ;
        RECT  2.140 1.760 2.400 2.555 ;
        RECT  1.630 0.405 2.240 0.585 ;
        RECT  1.950 1.760 2.140 1.920 ;
        RECT  0.955 2.395 2.140 2.555 ;
        RECT  1.790 0.855 1.950 1.920 ;
        RECT  1.520 0.355 1.630 0.585 ;
        RECT  1.360 0.355 1.520 2.210 ;
        RECT  1.000 0.690 1.160 2.075 ;
        RECT  0.930 0.690 1.000 0.975 ;
        RECT  0.915 1.685 1.000 2.075 ;
        RECT  0.695 2.305 0.955 2.555 ;
        RECT  0.125 0.815 0.930 0.975 ;
        RECT  0.605 1.685 0.915 1.945 ;
    END
END TBUFX4MTH

MACRO TBUFX6MTH
    CLASS CORE ;
    FOREIGN TBUFX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.510 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  4.125 0.445 4.410 2.455 ;
        RECT  3.185 0.445 4.125 0.715 ;
        RECT  3.160 2.095 4.125 2.365 ;
        END
        AntennaDiffArea 1.043 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 0.565 1.470 ;
        RECT  0.100 1.205 0.310 1.580 ;
        END
        AntennaGateArea 0.1508 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.360 1.280 2.770 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.935 -0.130 4.510 0.130 ;
        RECT  2.675 -0.130 2.935 0.715 ;
        RECT  0.810 -0.130 2.675 0.130 ;
        RECT  0.210 -0.130 0.810 0.485 ;
        RECT  0.000 -0.130 0.210 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.910 2.740 4.510 3.000 ;
        RECT  2.650 2.130 2.910 3.000 ;
        RECT  0.405 2.740 2.650 3.000 ;
        RECT  0.150 2.255 0.405 3.000 ;
        RECT  0.000 2.740 0.150 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.595 1.395 3.855 1.655 ;
        RECT  3.115 1.495 3.595 1.655 ;
        RECT  3.105 0.930 3.375 1.295 ;
        RECT  2.955 1.495 3.115 1.920 ;
        RECT  2.480 0.930 3.105 1.090 ;
        RECT  2.395 1.760 2.955 1.920 ;
        RECT  2.320 0.310 2.480 1.090 ;
        RECT  2.140 1.760 2.395 2.555 ;
        RECT  2.165 0.310 2.320 0.565 ;
        RECT  1.475 0.310 2.165 0.470 ;
        RECT  1.980 0.745 2.140 2.555 ;
        RECT  1.915 0.745 1.980 0.920 ;
        RECT  1.290 2.395 1.980 2.555 ;
        RECT  1.655 0.650 1.915 0.920 ;
        RECT  1.625 1.950 1.785 2.210 ;
        RECT  1.475 1.950 1.625 2.110 ;
        RECT  1.315 0.310 1.475 2.110 ;
        RECT  1.105 0.310 1.315 0.635 ;
        RECT  0.690 2.305 1.290 2.555 ;
        RECT  0.975 0.815 1.135 1.945 ;
        RECT  0.125 0.815 0.975 0.975 ;
        RECT  0.575 1.685 0.975 1.945 ;
    END
END TBUFX6MTH

MACRO TBUFX8MTH
    CLASS CORE ;
    FOREIGN TBUFX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.150 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT TRISTATE ;
        PORT
        LAYER METAL1 ;
        RECT  5.255 0.355 5.515 2.450 ;
        RECT  5.245 0.745 5.255 2.450 ;
        RECT  5.020 0.745 5.245 2.125 ;
        RECT  4.495 0.745 5.020 1.085 ;
        RECT  4.480 1.805 5.020 2.125 ;
        RECT  4.235 0.355 4.495 1.085 ;
        RECT  4.220 1.805 4.480 2.450 ;
        END
        AntennaDiffArea 1.131 ;
    END Y
    PIN OE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.080 0.505 1.680 ;
        END
        AntennaGateArea 0.2184 ;
    END OE
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.770 1.175 3.095 1.435 ;
        RECT  2.495 1.175 2.770 1.580 ;
        END
        AntennaGateArea 0.351 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.025 -0.130 6.150 0.130 ;
        RECT  5.765 -0.130 6.025 0.980 ;
        RECT  5.005 -0.130 5.765 0.130 ;
        RECT  4.745 -0.130 5.005 0.565 ;
        RECT  3.985 -0.130 4.745 0.130 ;
        RECT  3.725 -0.130 3.985 0.615 ;
        RECT  2.935 -0.130 3.725 0.130 ;
        RECT  2.675 -0.130 2.935 0.650 ;
        RECT  0.860 -0.130 2.675 0.130 ;
        RECT  0.260 -0.130 0.860 0.300 ;
        RECT  0.000 -0.130 0.260 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.020 2.740 6.150 3.000 ;
        RECT  5.760 1.815 6.020 3.000 ;
        RECT  4.995 2.740 5.760 3.000 ;
        RECT  4.735 2.305 4.995 3.000 ;
        RECT  3.970 2.740 4.735 3.000 ;
        RECT  3.710 1.890 3.970 3.000 ;
        RECT  2.925 2.740 3.710 3.000 ;
        RECT  2.665 2.160 2.925 3.000 ;
        RECT  0.535 2.740 2.665 3.000 ;
        RECT  0.275 2.570 0.535 3.000 ;
        RECT  0.000 2.740 0.275 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.275 1.435 4.535 1.625 ;
        RECT  3.455 1.465 4.275 1.625 ;
        RECT  3.950 1.125 4.050 1.285 ;
        RECT  3.790 0.830 3.950 1.285 ;
        RECT  3.470 0.830 3.790 0.995 ;
        RECT  3.210 0.590 3.470 0.995 ;
        RECT  3.295 1.465 3.455 2.360 ;
        RECT  3.195 1.760 3.295 2.360 ;
        RECT  2.375 0.830 3.210 0.995 ;
        RECT  2.365 1.760 3.195 1.920 ;
        RECT  2.215 0.310 2.375 0.995 ;
        RECT  2.270 1.760 2.365 2.220 ;
        RECT  2.110 1.305 2.270 2.220 ;
        RECT  1.405 0.310 2.215 0.470 ;
        RECT  1.915 1.305 2.110 1.465 ;
        RECT  1.325 2.060 2.110 2.220 ;
        RECT  1.755 0.655 1.915 1.465 ;
        RECT  1.615 1.645 1.875 1.880 ;
        RECT  0.880 2.400 1.875 2.560 ;
        RECT  1.655 0.655 1.755 0.915 ;
        RECT  1.405 1.645 1.615 1.805 ;
        RECT  1.245 0.310 1.405 1.805 ;
        RECT  1.065 2.030 1.325 2.220 ;
        RECT  1.145 0.540 1.245 0.800 ;
        RECT  0.880 0.985 1.065 1.245 ;
        RECT  0.720 0.700 0.880 2.560 ;
        RECT  0.415 0.700 0.720 0.860 ;
        RECT  0.175 1.880 0.720 2.140 ;
        RECT  0.155 0.600 0.415 0.860 ;
    END
END TBUFX8MTH

MACRO TIEHIMTH
    CLASS CORE ;
    FOREIGN TIEHIMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.000 1.700 1.130 1.990 ;
        RECT  0.740 1.700 1.000 2.390 ;
        END
        AntennaDiffArea 0.289 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 -0.130 1.230 0.130 ;
        RECT  0.200 -0.130 0.460 1.025 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 2.740 1.230 3.000 ;
        RECT  0.200 1.685 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.770 0.765 1.030 1.485 ;
        RECT  0.570 1.225 0.770 1.485 ;
    END
END TIEHIMTH

MACRO TIELOMTH
    CLASS CORE ;
    FOREIGN TIELOMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.230 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.740 0.425 1.130 1.025 ;
        END
        AntennaDiffArea 0.235 ;
    END Y
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 -0.130 1.230 0.130 ;
        RECT  0.200 -0.130 0.460 1.025 ;
        RECT  0.000 -0.130 0.200 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  0.460 2.740 1.230 3.000 ;
        RECT  0.200 1.690 0.460 3.000 ;
        RECT  0.000 2.740 0.200 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  0.780 1.225 1.040 1.945 ;
        RECT  0.570 1.225 0.780 1.485 ;
    END
END TIELOMTH

MACRO TLATNCAX12MTH
    CLASS CORE ;
    FOREIGN TLATNCAX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.940 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.425 0.810 13.225 2.005 ;
        RECT  11.805 0.810 12.425 1.145 ;
        RECT  11.040 0.810 11.805 2.035 ;
        RECT  9.835 0.810 11.040 1.145 ;
        RECT  9.230 0.810 9.835 2.100 ;
        END
        AntennaDiffArea 1.678 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.040 0.880 6.560 1.265 ;
        RECT  5.880 0.880 6.040 1.540 ;
        RECT  5.170 1.380 5.880 1.540 ;
        RECT  5.010 1.120 5.170 1.540 ;
        RECT  4.400 1.120 5.010 1.280 ;
        RECT  4.240 1.120 4.400 1.540 ;
        RECT  3.395 1.380 4.240 1.540 ;
        END
        AntennaGateArea 0.7865 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.410 1.225 1.080 1.580 ;
        END
        AntennaGateArea 0.5135 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.575 -0.130 13.940 0.130 ;
        RECT  13.315 -0.130 13.575 0.590 ;
        RECT  12.240 -0.130 13.315 0.130 ;
        RECT  11.300 -0.130 12.240 0.250 ;
        RECT  10.365 -0.130 11.300 0.130 ;
        RECT  10.105 -0.130 10.365 0.250 ;
        RECT  9.100 -0.130 10.105 0.130 ;
        RECT  8.840 -0.130 9.100 0.250 ;
        RECT  6.820 -0.130 8.840 0.130 ;
        RECT  6.560 -0.130 6.820 0.265 ;
        RECT  5.070 -0.130 6.560 0.130 ;
        RECT  4.810 -0.130 5.070 0.250 ;
        RECT  0.385 -0.130 4.810 0.130 ;
        RECT  0.125 -0.130 0.385 1.015 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.815 2.740 13.940 3.000 ;
        RECT  13.555 2.555 13.815 3.000 ;
        RECT  10.520 2.740 13.555 3.000 ;
        RECT  10.360 1.805 10.520 3.000 ;
        RECT  8.845 2.740 10.360 3.000 ;
        RECT  8.245 2.620 8.845 3.000 ;
        RECT  1.875 2.740 8.245 3.000 ;
        RECT  1.615 2.505 1.875 3.000 ;
        RECT  0.000 2.740 1.615 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  13.405 1.315 13.665 2.375 ;
        RECT  12.245 2.215 13.405 2.375 ;
        RECT  12.875 0.395 13.135 0.590 ;
        RECT  10.985 0.430 12.875 0.590 ;
        RECT  11.985 1.365 12.245 2.375 ;
        RECT  10.860 2.215 11.985 2.375 ;
        RECT  10.725 0.395 10.985 0.590 ;
        RECT  10.700 1.365 10.860 2.375 ;
        RECT  8.660 0.430 10.725 0.590 ;
        RECT  10.180 1.365 10.700 1.575 ;
        RECT  10.020 1.365 10.180 2.440 ;
        RECT  9.050 2.280 10.020 2.440 ;
        RECT  8.890 1.315 9.050 2.440 ;
        RECT  7.960 2.280 8.890 2.440 ;
        RECT  8.500 0.310 8.660 0.590 ;
        RECT  7.880 0.310 8.500 0.470 ;
        RECT  8.320 1.575 8.450 1.895 ;
        RECT  8.065 0.685 8.320 1.895 ;
        RECT  8.060 0.685 8.065 1.785 ;
        RECT  7.465 1.575 8.060 1.785 ;
        RECT  7.800 2.280 7.960 2.560 ;
        RECT  7.720 0.310 7.880 1.395 ;
        RECT  2.565 2.400 7.800 2.560 ;
        RECT  7.480 0.310 7.720 0.695 ;
        RECT  7.255 1.235 7.720 1.395 ;
        RECT  6.910 0.895 7.540 1.055 ;
        RECT  5.870 0.535 7.480 0.695 ;
        RECT  7.255 1.985 7.480 2.220 ;
        RECT  7.095 1.235 7.255 2.220 ;
        RECT  2.745 2.060 7.095 2.220 ;
        RECT  6.750 0.895 6.910 1.645 ;
        RECT  6.530 1.485 6.750 1.645 ;
        RECT  6.220 1.485 6.530 1.880 ;
        RECT  4.790 1.720 6.220 1.880 ;
        RECT  5.710 0.430 5.870 0.695 ;
        RECT  4.220 0.430 5.710 0.590 ;
        RECT  5.530 0.940 5.700 1.200 ;
        RECT  5.370 0.775 5.530 1.200 ;
        RECT  4.060 0.775 5.370 0.935 ;
        RECT  4.580 1.460 4.790 1.880 ;
        RECT  3.175 1.720 4.580 1.880 ;
        RECT  3.960 0.405 4.220 0.590 ;
        RECT  3.900 0.775 4.060 1.195 ;
        RECT  2.400 0.405 3.960 0.565 ;
        RECT  2.995 0.775 3.900 0.935 ;
        RECT  2.915 1.495 3.175 1.880 ;
        RECT  2.830 0.745 2.995 0.935 ;
        RECT  2.450 1.720 2.915 1.880 ;
        RECT  2.570 0.745 2.830 1.145 ;
        RECT  2.220 0.745 2.570 0.905 ;
        RECT  2.405 2.165 2.565 2.560 ;
        RECT  2.315 1.720 2.450 1.985 ;
        RECT  1.485 2.165 2.405 2.325 ;
        RECT  2.155 1.105 2.315 1.985 ;
        RECT  2.060 0.395 2.220 0.905 ;
        RECT  1.880 1.105 2.155 1.265 ;
        RECT  1.485 0.395 2.060 0.555 ;
        RECT  1.485 1.445 1.975 1.605 ;
        RECT  1.720 0.765 1.880 1.265 ;
        RECT  1.325 0.395 1.485 2.380 ;
        RECT  0.925 0.395 1.325 0.555 ;
        RECT  1.065 1.780 1.325 2.380 ;
        RECT  0.385 1.780 1.065 2.000 ;
        RECT  0.665 0.395 0.925 0.995 ;
        RECT  0.125 1.780 0.385 2.380 ;
    END
END TLATNCAX12MTH

MACRO TLATNCAX16MTH
    CLASS CORE ;
    FOREIGN TLATNCAX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 15.580 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  14.245 0.810 15.005 2.020 ;
        RECT  13.005 0.810 14.245 1.185 ;
        RECT  12.465 0.810 13.005 2.035 ;
        RECT  11.765 0.810 12.465 1.185 ;
        RECT  11.080 0.810 11.765 2.035 ;
        RECT  9.800 0.810 11.080 1.185 ;
        RECT  9.230 0.810 9.800 2.100 ;
        END
        AntennaDiffArea 2.262 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.040 0.880 6.560 1.265 ;
        RECT  5.880 0.880 6.040 1.540 ;
        RECT  5.170 1.380 5.880 1.540 ;
        RECT  5.010 1.110 5.170 1.540 ;
        RECT  4.400 1.110 5.010 1.270 ;
        RECT  4.240 1.110 4.400 1.540 ;
        RECT  3.395 1.380 4.240 1.540 ;
        END
        AntennaGateArea 0.7865 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.410 1.225 1.080 1.580 ;
        END
        AntennaGateArea 0.5161 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.405 -0.130 15.580 0.130 ;
        RECT  15.245 -0.130 15.405 1.000 ;
        RECT  14.235 -0.130 15.245 0.130 ;
        RECT  13.295 -0.130 14.235 0.250 ;
        RECT  12.170 -0.130 13.295 0.130 ;
        RECT  11.230 -0.130 12.170 0.250 ;
        RECT  10.365 -0.130 11.230 0.130 ;
        RECT  10.105 -0.130 10.365 0.250 ;
        RECT  9.100 -0.130 10.105 0.130 ;
        RECT  8.840 -0.130 9.100 0.250 ;
        RECT  6.810 -0.130 8.840 0.130 ;
        RECT  6.550 -0.130 6.810 0.355 ;
        RECT  5.070 -0.130 6.550 0.130 ;
        RECT  4.810 -0.130 5.070 0.250 ;
        RECT  0.385 -0.130 4.810 0.130 ;
        RECT  0.125 -0.130 0.385 1.015 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.455 2.740 15.580 3.000 ;
        RECT  15.195 2.570 15.455 3.000 ;
        RECT  13.725 2.740 15.195 3.000 ;
        RECT  13.565 1.810 13.725 3.000 ;
        RECT  10.520 2.740 13.565 3.000 ;
        RECT  10.360 1.805 10.520 3.000 ;
        RECT  8.845 2.740 10.360 3.000 ;
        RECT  8.245 2.620 8.845 3.000 ;
        RECT  1.875 2.740 8.245 3.000 ;
        RECT  1.615 2.505 1.875 3.000 ;
        RECT  0.000 2.740 1.615 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.210 1.315 15.370 2.390 ;
        RECT  14.065 2.230 15.210 2.390 ;
        RECT  14.465 0.400 14.725 0.590 ;
        RECT  13.045 0.430 14.465 0.590 ;
        RECT  13.905 1.365 14.065 2.390 ;
        RECT  13.385 1.365 13.905 1.575 ;
        RECT  13.225 1.365 13.385 2.375 ;
        RECT  12.245 2.215 13.225 2.375 ;
        RECT  12.785 0.400 13.045 0.590 ;
        RECT  10.985 0.430 12.785 0.590 ;
        RECT  11.985 1.365 12.245 2.375 ;
        RECT  10.860 2.215 11.985 2.375 ;
        RECT  10.725 0.400 10.985 0.590 ;
        RECT  10.700 1.365 10.860 2.375 ;
        RECT  8.660 0.430 10.725 0.590 ;
        RECT  10.180 1.365 10.700 1.575 ;
        RECT  10.020 1.365 10.180 2.440 ;
        RECT  9.050 2.280 10.020 2.440 ;
        RECT  8.890 1.315 9.050 2.440 ;
        RECT  7.960 2.280 8.890 2.440 ;
        RECT  8.500 0.310 8.660 0.590 ;
        RECT  7.880 0.310 8.500 0.470 ;
        RECT  8.320 1.575 8.450 1.895 ;
        RECT  8.065 0.685 8.320 1.895 ;
        RECT  8.060 0.685 8.065 1.785 ;
        RECT  7.465 1.575 8.060 1.785 ;
        RECT  7.800 2.280 7.960 2.560 ;
        RECT  7.720 0.310 7.880 1.395 ;
        RECT  2.565 2.400 7.800 2.560 ;
        RECT  7.480 0.310 7.720 0.695 ;
        RECT  7.255 1.235 7.720 1.395 ;
        RECT  6.910 0.895 7.540 1.055 ;
        RECT  5.870 0.535 7.480 0.695 ;
        RECT  7.255 2.030 7.480 2.220 ;
        RECT  7.095 1.235 7.255 2.220 ;
        RECT  2.745 2.060 7.095 2.220 ;
        RECT  6.750 0.895 6.910 1.645 ;
        RECT  6.530 1.485 6.750 1.645 ;
        RECT  6.220 1.485 6.530 1.880 ;
        RECT  4.790 1.720 6.220 1.880 ;
        RECT  5.710 0.430 5.870 0.695 ;
        RECT  3.405 0.430 5.710 0.590 ;
        RECT  5.530 0.940 5.700 1.200 ;
        RECT  5.370 0.770 5.530 1.200 ;
        RECT  4.060 0.770 5.370 0.930 ;
        RECT  4.580 1.460 4.790 1.880 ;
        RECT  3.175 1.720 4.580 1.880 ;
        RECT  3.900 0.770 4.060 1.195 ;
        RECT  2.830 0.770 3.900 0.930 ;
        RECT  3.245 0.405 3.405 0.590 ;
        RECT  2.400 0.405 3.245 0.565 ;
        RECT  2.915 1.495 3.175 1.880 ;
        RECT  2.490 1.720 2.915 1.880 ;
        RECT  2.730 0.770 2.830 1.145 ;
        RECT  2.570 0.745 2.730 1.145 ;
        RECT  2.220 0.745 2.570 0.905 ;
        RECT  2.405 2.165 2.565 2.560 ;
        RECT  2.315 1.720 2.490 1.985 ;
        RECT  1.485 2.165 2.405 2.325 ;
        RECT  2.155 1.085 2.315 1.985 ;
        RECT  2.060 0.395 2.220 0.905 ;
        RECT  1.880 1.085 2.155 1.245 ;
        RECT  1.485 0.395 2.060 0.555 ;
        RECT  1.485 1.425 1.975 1.585 ;
        RECT  1.720 0.765 1.880 1.245 ;
        RECT  1.325 0.395 1.485 2.380 ;
        RECT  0.925 0.395 1.325 0.555 ;
        RECT  1.065 1.780 1.325 2.380 ;
        RECT  0.385 1.780 1.065 2.000 ;
        RECT  0.665 0.395 0.925 0.995 ;
        RECT  0.125 1.780 0.385 2.380 ;
    END
END TLATNCAX16MTH

MACRO TLATNCAX20MTH
    CLASS CORE ;
    FOREIGN TLATNCAX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 20.090 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  18.755 0.810 19.510 2.045 ;
        RECT  17.860 0.810 18.755 1.185 ;
        RECT  17.265 0.810 17.860 1.995 ;
        RECT  16.065 0.810 17.265 1.185 ;
        RECT  15.465 0.810 16.065 2.035 ;
        RECT  14.840 0.810 15.465 1.185 ;
        RECT  14.125 0.810 14.840 2.035 ;
        RECT  12.820 0.810 14.125 1.185 ;
        RECT  12.265 0.810 12.820 2.100 ;
        END
        AntennaDiffArea 2.898 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 0.880 9.595 1.265 ;
        RECT  8.915 0.880 9.075 1.540 ;
        RECT  8.205 1.380 8.915 1.540 ;
        RECT  8.045 1.110 8.205 1.540 ;
        RECT  7.435 1.110 8.045 1.270 ;
        RECT  7.275 1.110 7.435 1.540 ;
        RECT  6.640 1.380 7.275 1.540 ;
        RECT  6.430 1.260 6.640 1.540 ;
        RECT  4.680 1.260 6.430 1.420 ;
        END
        AntennaGateArea 1.0166 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.440 1.225 2.085 1.580 ;
        END
        AntennaGateArea 1.0192 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  19.865 -0.130 20.090 0.130 ;
        RECT  18.925 -0.130 19.865 0.300 ;
        RECT  18.195 -0.130 18.925 0.130 ;
        RECT  17.935 -0.130 18.195 0.250 ;
        RECT  17.025 -0.130 17.935 0.130 ;
        RECT  16.085 -0.130 17.025 0.250 ;
        RECT  15.135 -0.130 16.085 0.130 ;
        RECT  14.195 -0.130 15.135 0.250 ;
        RECT  13.400 -0.130 14.195 0.130 ;
        RECT  13.140 -0.130 13.400 0.250 ;
        RECT  12.135 -0.130 13.140 0.130 ;
        RECT  11.875 -0.130 12.135 0.250 ;
        RECT  9.855 -0.130 11.875 0.130 ;
        RECT  9.595 -0.130 9.855 0.265 ;
        RECT  8.105 -0.130 9.595 0.130 ;
        RECT  7.845 -0.130 8.105 0.250 ;
        RECT  4.845 -0.130 7.845 0.130 ;
        RECT  4.585 -0.130 4.845 0.250 ;
        RECT  1.825 -0.130 4.585 0.130 ;
        RECT  1.565 -0.130 1.825 0.615 ;
        RECT  0.000 -0.130 1.565 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.745 2.740 20.090 3.000 ;
        RECT  16.585 1.915 16.745 3.000 ;
        RECT  13.605 2.740 16.585 3.000 ;
        RECT  13.345 1.805 13.605 3.000 ;
        RECT  11.880 2.740 13.345 3.000 ;
        RECT  11.280 2.620 11.880 3.000 ;
        RECT  5.140 2.740 11.280 3.000 ;
        RECT  4.880 2.620 5.140 3.000 ;
        RECT  3.135 2.740 4.880 3.000 ;
        RECT  2.875 2.505 3.135 3.000 ;
        RECT  1.915 2.740 2.875 3.000 ;
        RECT  1.655 2.160 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.160 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  19.725 1.295 19.885 2.425 ;
        RECT  18.300 2.265 19.725 2.425 ;
        RECT  18.480 0.395 18.740 0.590 ;
        RECT  17.760 0.430 18.480 0.590 ;
        RECT  18.040 1.365 18.300 2.425 ;
        RECT  17.085 2.265 18.040 2.425 ;
        RECT  17.160 0.395 17.760 0.590 ;
        RECT  15.900 0.430 17.160 0.590 ;
        RECT  16.925 1.365 17.085 2.425 ;
        RECT  16.405 1.365 16.925 1.575 ;
        RECT  16.245 1.365 16.405 2.375 ;
        RECT  15.280 2.215 16.245 2.375 ;
        RECT  15.640 0.395 15.900 0.590 ;
        RECT  14.020 0.430 15.640 0.590 ;
        RECT  15.020 1.365 15.280 2.375 ;
        RECT  13.945 2.215 15.020 2.375 ;
        RECT  13.760 0.395 14.020 0.590 ;
        RECT  13.785 1.365 13.945 2.375 ;
        RECT  13.160 1.365 13.785 1.575 ;
        RECT  11.695 0.430 13.760 0.590 ;
        RECT  13.000 1.365 13.160 2.440 ;
        RECT  12.085 2.280 13.000 2.440 ;
        RECT  11.925 1.315 12.085 2.440 ;
        RECT  10.995 2.280 11.925 2.440 ;
        RECT  11.535 0.310 11.695 0.590 ;
        RECT  10.915 0.310 11.535 0.470 ;
        RECT  11.355 1.575 11.485 1.895 ;
        RECT  11.100 0.685 11.355 1.895 ;
        RECT  11.095 0.685 11.100 1.785 ;
        RECT  10.500 1.575 11.095 1.785 ;
        RECT  10.835 2.280 10.995 2.560 ;
        RECT  10.755 0.310 10.915 1.395 ;
        RECT  5.480 2.400 10.835 2.560 ;
        RECT  10.515 0.310 10.755 0.695 ;
        RECT  10.290 1.235 10.755 1.395 ;
        RECT  9.945 0.895 10.575 1.055 ;
        RECT  8.905 0.535 10.515 0.695 ;
        RECT  10.290 1.985 10.515 2.220 ;
        RECT  10.130 1.235 10.290 2.220 ;
        RECT  5.820 2.060 10.130 2.220 ;
        RECT  9.785 0.895 9.945 1.645 ;
        RECT  9.565 1.485 9.785 1.645 ;
        RECT  9.255 1.485 9.565 1.880 ;
        RECT  7.825 1.720 9.255 1.880 ;
        RECT  8.745 0.430 8.905 0.695 ;
        RECT  4.480 0.430 8.745 0.590 ;
        RECT  8.565 0.940 8.735 1.200 ;
        RECT  8.405 0.770 8.565 1.200 ;
        RECT  7.095 0.770 8.405 0.930 ;
        RECT  7.615 1.465 7.825 1.880 ;
        RECT  6.195 1.720 7.615 1.880 ;
        RECT  6.935 0.770 7.095 1.195 ;
        RECT  5.865 0.770 6.935 0.930 ;
        RECT  6.000 1.600 6.195 1.880 ;
        RECT  3.780 1.600 6.000 1.760 ;
        RECT  5.605 0.770 5.865 1.080 ;
        RECT  5.660 1.940 5.820 2.220 ;
        RECT  4.290 1.940 5.660 2.100 ;
        RECT  4.165 0.770 5.605 0.930 ;
        RECT  5.320 2.280 5.480 2.560 ;
        RECT  4.700 2.280 5.320 2.440 ;
        RECT  4.540 2.280 4.700 2.555 ;
        RECT  3.670 2.395 4.540 2.555 ;
        RECT  4.320 0.405 4.480 0.590 ;
        RECT  3.735 0.405 4.320 0.565 ;
        RECT  4.030 1.940 4.290 2.215 ;
        RECT  4.095 0.770 4.165 1.075 ;
        RECT  3.905 0.745 4.095 1.075 ;
        RECT  3.555 0.745 3.905 0.905 ;
        RECT  3.645 1.600 3.780 1.985 ;
        RECT  3.510 2.165 3.670 2.555 ;
        RECT  3.485 1.085 3.645 1.985 ;
        RECT  3.395 0.395 3.555 0.905 ;
        RECT  2.495 2.165 3.510 2.325 ;
        RECT  3.215 1.085 3.485 1.245 ;
        RECT  2.495 0.395 3.395 0.555 ;
        RECT  2.495 1.425 3.305 1.585 ;
        RECT  3.055 0.765 3.215 1.245 ;
        RECT  2.335 0.395 2.495 2.405 ;
        RECT  2.075 0.395 2.335 0.995 ;
        RECT  2.235 1.805 2.335 2.405 ;
        RECT  1.405 1.805 2.235 1.980 ;
        RECT  1.315 0.835 2.075 0.995 ;
        RECT  1.145 1.805 1.405 2.410 ;
        RECT  1.055 0.395 1.315 0.995 ;
        RECT  0.385 1.805 1.145 1.980 ;
        RECT  0.385 0.835 1.055 0.995 ;
        RECT  0.125 0.395 0.385 0.995 ;
        RECT  0.125 1.805 0.385 2.405 ;
    END
END TLATNCAX20MTH

MACRO TLATNCAX2MTH
    CLASS CORE ;
    FOREIGN TLATNCAX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.330 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.070 0.770 5.230 2.415 ;
        RECT  4.540 0.770 5.070 0.930 ;
        RECT  4.900 1.700 5.070 2.415 ;
        END
        AntennaDiffArea 0.416 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.475 0.880 1.950 1.285 ;
        END
        AntennaGateArea 0.1729 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.055 0.355 2.025 ;
        END
        AntennaGateArea 0.1378 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.260 -0.130 5.330 0.130 ;
        RECT  3.320 -0.130 4.260 0.250 ;
        RECT  0.385 -0.130 3.320 0.130 ;
        RECT  0.125 -0.130 0.385 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.210 2.740 5.330 3.000 ;
        RECT  3.270 2.570 4.210 3.000 ;
        RECT  1.525 2.740 3.270 3.000 ;
        RECT  1.265 2.515 1.525 3.000 ;
        RECT  0.000 2.740 1.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.715 0.390 4.975 0.590 ;
        RECT  3.115 0.430 4.715 0.590 ;
        RECT  4.250 1.250 4.510 2.360 ;
        RECT  3.005 2.200 4.250 2.360 ;
        RECT  3.745 0.770 3.905 1.945 ;
        RECT  3.565 0.770 3.745 0.975 ;
        RECT  2.995 1.680 3.745 1.945 ;
        RECT  2.635 1.250 3.565 1.410 ;
        RECT  2.955 0.430 3.115 0.845 ;
        RECT  2.845 2.200 3.005 2.560 ;
        RECT  2.635 0.685 2.955 0.845 ;
        RECT  1.865 2.400 2.845 2.560 ;
        RECT  1.225 0.310 2.775 0.470 ;
        RECT  2.475 0.685 2.635 2.190 ;
        RECT  2.245 0.685 2.475 0.845 ;
        RECT  2.205 2.030 2.475 2.190 ;
        RECT  2.135 1.025 2.295 1.765 ;
        RECT  1.865 1.605 2.135 1.765 ;
        RECT  1.705 1.605 1.865 2.560 ;
        RECT  0.775 2.175 1.705 2.335 ;
        RECT  1.065 0.310 1.225 1.970 ;
        RECT  0.965 0.310 1.065 0.565 ;
        RECT  0.925 1.710 1.065 1.970 ;
        RECT  0.735 1.270 0.885 1.530 ;
        RECT  0.695 2.175 0.775 2.470 ;
        RECT  0.695 0.765 0.735 1.530 ;
        RECT  0.535 0.765 0.695 2.470 ;
    END
END TLATNCAX2MTH

MACRO TLATNCAX3MTH
    CLASS CORE ;
    FOREIGN TLATNCAX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.815 0.420 5.075 2.085 ;
        RECT  4.610 1.645 4.815 2.085 ;
        END
        AntennaDiffArea 0.428 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.555 0.880 1.965 1.380 ;
        END
        AntennaGateArea 0.1885 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.355 2.135 ;
        END
        AntennaGateArea 0.1846 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.615 -0.130 5.740 0.130 ;
        RECT  5.355 -0.130 5.615 0.775 ;
        RECT  4.525 -0.130 5.355 0.130 ;
        RECT  4.265 -0.130 4.525 0.775 ;
        RECT  3.445 -0.130 4.265 0.130 ;
        RECT  3.185 -0.130 3.445 0.335 ;
        RECT  0.385 -0.130 3.185 0.130 ;
        RECT  0.125 -0.130 0.385 1.025 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.925 2.740 5.740 3.000 ;
        RECT  3.325 2.600 3.925 3.000 ;
        RECT  1.525 2.740 3.325 3.000 ;
        RECT  1.265 2.560 1.525 3.000 ;
        RECT  0.000 2.740 1.265 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.445 1.045 5.545 1.645 ;
        RECT  5.285 1.045 5.445 2.480 ;
        RECT  4.355 2.320 5.285 2.480 ;
        RECT  4.195 1.195 4.355 2.480 ;
        RECT  3.145 2.255 4.195 2.415 ;
        RECT  3.855 0.515 4.015 1.940 ;
        RECT  3.695 0.515 3.855 0.775 ;
        RECT  2.985 1.590 3.855 1.940 ;
        RECT  2.785 1.010 3.675 1.270 ;
        RECT  2.985 2.255 3.145 2.560 ;
        RECT  1.865 2.400 2.985 2.560 ;
        RECT  1.335 0.310 2.875 0.470 ;
        RECT  2.625 0.680 2.785 2.190 ;
        RECT  2.355 0.680 2.625 0.840 ;
        RECT  2.205 2.030 2.625 2.190 ;
        RECT  2.345 1.055 2.445 1.215 ;
        RECT  2.185 1.055 2.345 1.765 ;
        RECT  1.865 1.605 2.185 1.765 ;
        RECT  1.705 1.605 1.865 2.560 ;
        RECT  0.805 2.210 1.705 2.370 ;
        RECT  1.175 0.310 1.335 1.945 ;
        RECT  1.075 0.310 1.175 0.565 ;
        RECT  0.925 1.685 1.175 1.945 ;
        RECT  0.725 0.765 0.985 1.495 ;
        RECT  0.725 2.210 0.805 2.470 ;
        RECT  0.565 0.765 0.725 2.470 ;
    END
END TLATNCAX3MTH

MACRO TLATNCAX4MTH
    CLASS CORE ;
    FOREIGN TLATNCAX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.070 0.505 7.280 2.125 ;
        RECT  5.840 0.505 7.070 0.785 ;
        RECT  6.410 1.865 7.070 2.125 ;
        RECT  6.150 1.865 6.410 2.465 ;
        END
        AntennaDiffArea 0.572 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.950 1.235 3.145 1.495 ;
        RECT  1.630 1.235 1.950 1.580 ;
        END
        AntennaGateArea 0.2652 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.155 0.540 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.015 -0.130 7.380 0.130 ;
        RECT  6.415 -0.130 7.015 0.315 ;
        RECT  3.735 -0.130 6.415 0.130 ;
        RECT  3.135 -0.130 3.735 0.250 ;
        RECT  1.655 -0.130 3.135 0.130 ;
        RECT  0.715 -0.130 1.655 0.250 ;
        RECT  0.000 -0.130 0.715 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.230 2.740 7.380 3.000 ;
        RECT  6.970 2.305 7.230 3.000 ;
        RECT  5.500 2.740 6.970 3.000 ;
        RECT  5.000 2.195 5.500 3.000 ;
        RECT  1.670 2.740 5.000 3.000 ;
        RECT  0.730 2.610 1.670 3.000 ;
        RECT  0.000 2.740 0.730 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.680 1.000 6.840 1.260 ;
        RECT  5.760 1.000 6.680 1.160 ;
        RECT  5.980 1.365 6.240 1.685 ;
        RECT  5.275 1.525 5.980 1.685 ;
        RECT  5.655 1.000 5.760 1.325 ;
        RECT  5.495 0.310 5.655 1.325 ;
        RECT  4.110 0.310 5.495 0.470 ;
        RECT  5.115 0.650 5.275 1.945 ;
        RECT  4.445 0.650 5.115 0.810 ;
        RECT  4.975 1.685 5.115 1.945 ;
        RECT  4.785 1.005 4.935 1.265 ;
        RECT  4.625 1.005 4.785 2.560 ;
        RECT  2.710 2.400 4.625 2.560 ;
        RECT  4.285 0.650 4.445 2.220 ;
        RECT  3.485 2.060 4.285 2.220 ;
        RECT  3.950 0.310 4.110 0.590 ;
        RECT  3.920 0.770 4.105 1.880 ;
        RECT  2.715 0.430 3.950 0.590 ;
        RECT  3.665 0.770 3.920 0.930 ;
        RECT  3.665 1.720 3.920 1.880 ;
        RECT  3.485 1.215 3.625 1.475 ;
        RECT  3.325 0.810 3.485 2.220 ;
        RECT  2.285 0.810 3.325 0.970 ;
        RECT  2.545 1.755 3.325 1.915 ;
        RECT  2.115 0.310 2.715 0.590 ;
        RECT  2.115 2.270 2.710 2.560 ;
        RECT  2.285 1.755 2.545 2.090 ;
        RECT  0.880 0.430 2.115 0.590 ;
        RECT  1.345 2.270 2.115 2.430 ;
        RECT  1.185 0.815 1.345 2.430 ;
        RECT  1.065 0.815 1.185 0.975 ;
        RECT  1.065 1.695 1.185 2.430 ;
        RECT  0.880 1.245 0.995 1.505 ;
        RECT  0.720 0.430 0.880 1.965 ;
        RECT  0.385 0.815 0.720 0.975 ;
        RECT  0.385 1.805 0.720 1.965 ;
        RECT  0.125 0.375 0.385 0.975 ;
        RECT  0.125 1.805 0.385 2.405 ;
    END
END TLATNCAX4MTH

MACRO TLATNCAX6MTH
    CLASS CORE ;
    FOREIGN TLATNCAX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.225 0.770 8.510 2.400 ;
        RECT  6.845 0.770 8.225 1.040 ;
        RECT  6.575 0.770 6.845 2.100 ;
        END
        AntennaDiffArea 1.048 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.135 0.880 3.615 1.265 ;
        RECT  2.975 0.880 3.135 1.540 ;
        RECT  2.125 1.380 2.975 1.540 ;
        END
        AntennaGateArea 0.3016 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.135 0.565 1.735 ;
        END
        AntennaGateArea 0.3289 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.480 -0.130 8.610 0.130 ;
        RECT  8.220 -0.130 8.480 0.590 ;
        RECT  7.460 -0.130 8.220 0.130 ;
        RECT  7.200 -0.130 7.460 0.250 ;
        RECT  6.195 -0.130 7.200 0.130 ;
        RECT  5.935 -0.130 6.195 0.250 ;
        RECT  3.905 -0.130 5.935 0.130 ;
        RECT  3.645 -0.130 3.905 0.250 ;
        RECT  2.085 -0.130 3.645 0.130 ;
        RECT  1.145 -0.130 2.085 0.250 ;
        RECT  0.000 -0.130 1.145 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.665 2.740 8.610 3.000 ;
        RECT  7.405 1.805 7.665 3.000 ;
        RECT  5.940 2.740 7.405 3.000 ;
        RECT  5.340 2.620 5.940 3.000 ;
        RECT  2.295 2.740 5.340 3.000 ;
        RECT  1.355 2.620 2.295 3.000 ;
        RECT  0.000 2.740 1.355 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.780 0.395 8.040 0.590 ;
        RECT  5.755 0.430 7.780 0.590 ;
        RECT  7.185 1.315 7.495 1.575 ;
        RECT  7.025 1.315 7.185 2.440 ;
        RECT  6.195 2.280 7.025 2.440 ;
        RECT  5.935 1.365 6.195 2.440 ;
        RECT  5.055 2.280 5.935 2.440 ;
        RECT  5.595 0.310 5.755 0.590 ;
        RECT  4.975 0.310 5.595 0.470 ;
        RECT  5.415 1.450 5.545 1.895 ;
        RECT  5.285 0.685 5.415 1.895 ;
        RECT  5.155 0.685 5.285 1.730 ;
        RECT  4.575 1.450 5.155 1.730 ;
        RECT  4.895 2.280 5.055 2.560 ;
        RECT  4.815 0.310 4.975 1.270 ;
        RECT  2.860 2.400 4.895 2.560 ;
        RECT  4.575 0.310 4.815 0.590 ;
        RECT  4.330 1.110 4.815 1.270 ;
        RECT  3.955 0.770 4.635 0.930 ;
        RECT  2.965 0.430 4.575 0.590 ;
        RECT  4.330 2.030 4.575 2.220 ;
        RECT  4.170 1.110 4.330 2.220 ;
        RECT  3.070 2.060 4.170 2.220 ;
        RECT  3.795 0.770 3.955 1.645 ;
        RECT  3.575 1.485 3.795 1.645 ;
        RECT  3.315 1.485 3.575 1.880 ;
        RECT  1.850 1.720 3.315 1.880 ;
        RECT  2.805 0.430 2.965 0.690 ;
        RECT  2.700 2.280 2.860 2.560 ;
        RECT  2.625 0.940 2.795 1.200 ;
        RECT  0.905 2.280 2.700 2.440 ;
        RECT  2.465 0.430 2.625 1.200 ;
        RECT  0.905 0.430 2.465 0.590 ;
        RECT  1.690 0.770 1.850 2.100 ;
        RECT  1.445 0.770 1.690 0.930 ;
        RECT  1.475 1.720 1.690 2.100 ;
        RECT  0.905 1.215 1.510 1.475 ;
        RECT  0.785 0.430 0.905 2.440 ;
        RECT  0.745 0.430 0.785 2.515 ;
        RECT  0.525 0.430 0.745 0.700 ;
        RECT  0.525 1.915 0.745 2.515 ;
    END
END TLATNCAX6MTH

MACRO TLATNCAX8MTH
    CLASS CORE ;
    FOREIGN TLATNCAX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.550 0.770 8.905 1.065 ;
        RECT  8.190 0.770 8.550 2.150 ;
        RECT  6.845 0.770 8.190 1.065 ;
        RECT  6.525 0.770 6.845 2.100 ;
        END
        AntennaDiffArea 1.214 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.135 0.880 3.615 1.265 ;
        RECT  2.975 0.880 3.135 1.540 ;
        RECT  2.125 1.380 2.975 1.540 ;
        END
        AntennaGateArea 0.3016 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.360 1.220 0.925 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.215 -0.130 9.430 0.130 ;
        RECT  8.275 -0.130 9.215 0.420 ;
        RECT  7.460 -0.130 8.275 0.130 ;
        RECT  7.200 -0.130 7.460 0.250 ;
        RECT  6.195 -0.130 7.200 0.130 ;
        RECT  5.935 -0.130 6.195 0.250 ;
        RECT  3.910 -0.130 5.935 0.130 ;
        RECT  3.650 -0.130 3.910 0.335 ;
        RECT  2.100 -0.130 3.650 0.130 ;
        RECT  1.160 -0.130 2.100 0.250 ;
        RECT  0.000 -0.130 1.160 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.255 2.740 9.430 3.000 ;
        RECT  9.095 1.825 9.255 3.000 ;
        RECT  7.665 2.740 9.095 3.000 ;
        RECT  7.405 1.805 7.665 3.000 ;
        RECT  5.940 2.740 7.405 3.000 ;
        RECT  5.340 2.620 5.940 3.000 ;
        RECT  2.480 2.740 5.340 3.000 ;
        RECT  1.540 2.620 2.480 3.000 ;
        RECT  1.330 2.740 1.540 3.000 ;
        RECT  1.070 2.620 1.330 3.000 ;
        RECT  0.000 2.740 1.070 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.915 1.245 9.135 1.505 ;
        RECT  8.755 1.245 8.915 2.490 ;
        RECT  8.005 2.330 8.755 2.490 ;
        RECT  7.820 0.310 8.080 0.590 ;
        RECT  7.845 1.315 8.005 2.490 ;
        RECT  7.185 1.315 7.845 1.575 ;
        RECT  5.755 0.430 7.820 0.590 ;
        RECT  7.025 1.315 7.185 2.440 ;
        RECT  6.195 2.280 7.025 2.440 ;
        RECT  5.935 1.365 6.195 2.440 ;
        RECT  5.055 2.280 5.935 2.440 ;
        RECT  5.595 0.310 5.755 0.590 ;
        RECT  4.975 0.310 5.595 0.470 ;
        RECT  5.415 1.530 5.545 1.895 ;
        RECT  5.280 0.705 5.415 1.895 ;
        RECT  5.155 0.705 5.280 1.795 ;
        RECT  4.575 1.535 5.155 1.795 ;
        RECT  4.895 2.280 5.055 2.560 ;
        RECT  4.815 0.310 4.975 1.355 ;
        RECT  2.860 2.400 4.895 2.560 ;
        RECT  4.575 0.310 4.815 0.675 ;
        RECT  4.330 1.195 4.815 1.355 ;
        RECT  3.955 0.855 4.635 1.015 ;
        RECT  2.965 0.515 4.575 0.675 ;
        RECT  4.330 2.030 4.575 2.220 ;
        RECT  4.170 1.195 4.330 2.220 ;
        RECT  3.070 2.060 4.170 2.220 ;
        RECT  3.795 0.855 3.955 1.645 ;
        RECT  3.625 1.485 3.795 1.645 ;
        RECT  3.315 1.485 3.625 1.880 ;
        RECT  1.850 1.720 3.315 1.880 ;
        RECT  2.805 0.415 2.965 0.675 ;
        RECT  2.700 2.280 2.860 2.560 ;
        RECT  2.625 0.940 2.795 1.200 ;
        RECT  1.265 2.280 2.700 2.440 ;
        RECT  2.465 0.430 2.625 1.200 ;
        RECT  1.265 0.430 2.465 0.590 ;
        RECT  1.690 0.770 1.850 2.100 ;
        RECT  1.445 0.770 1.690 0.930 ;
        RECT  1.475 1.720 1.690 2.100 ;
        RECT  1.265 1.215 1.510 1.475 ;
        RECT  1.105 0.430 1.265 2.440 ;
        RECT  0.785 0.430 1.105 0.590 ;
        RECT  0.785 2.280 1.105 2.440 ;
        RECT  0.525 0.430 0.785 0.930 ;
        RECT  0.525 1.840 0.785 2.440 ;
    END
END TLATNCAX8MTH

MACRO TLATNSRX1MTH
    CLASS CORE ;
    FOREIGN TLATNSRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.020 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.165 0.445 1.580 ;
        END
        AntennaGateArea 0.1157 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.855 0.315 3.955 0.475 ;
        RECT  3.695 0.315 3.855 1.140 ;
        RECT  2.865 0.980 3.695 1.140 ;
        RECT  2.705 0.685 2.865 1.220 ;
        RECT  1.950 0.685 2.705 0.845 ;
        RECT  1.790 0.685 1.950 1.580 ;
        RECT  1.740 1.150 1.790 1.580 ;
        END
        AntennaGateArea 0.1872 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.685 0.755 8.920 2.075 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.875 1.290 8.135 1.580 ;
        RECT  7.615 0.815 7.875 2.070 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  6.640 0.880 6.910 1.130 ;
        RECT  6.475 0.880 6.640 1.370 ;
        RECT  6.365 1.110 6.475 1.370 ;
        END
        AntennaGateArea 0.0754 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.025 2.435 1.580 ;
        END
        AntennaGateArea 0.1521 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.355 -0.130 9.020 0.130 ;
        RECT  7.415 -0.130 8.355 0.250 ;
        RECT  7.155 -0.130 7.415 0.130 ;
        RECT  6.215 -0.130 7.155 0.250 ;
        RECT  5.955 -0.130 6.215 0.130 ;
        RECT  5.015 -0.130 5.955 0.250 ;
        RECT  1.220 -0.130 5.015 0.130 ;
        RECT  0.280 -0.130 1.220 0.330 ;
        RECT  0.000 -0.130 0.280 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.385 2.740 9.020 3.000 ;
        RECT  8.125 1.815 8.385 3.000 ;
        RECT  7.625 2.740 8.125 3.000 ;
        RECT  6.685 2.555 7.625 3.000 ;
        RECT  5.165 2.740 6.685 3.000 ;
        RECT  4.665 2.185 5.165 3.000 ;
        RECT  2.065 2.740 4.665 3.000 ;
        RECT  1.465 2.520 2.065 3.000 ;
        RECT  0.725 2.740 1.465 3.000 ;
        RECT  0.125 2.465 0.725 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.345 0.430 8.505 1.485 ;
        RECT  7.365 0.430 8.345 0.590 ;
        RECT  7.205 0.430 7.365 2.025 ;
        RECT  7.105 0.430 7.205 0.960 ;
        RECT  7.105 1.865 7.205 2.025 ;
        RECT  5.015 0.430 7.105 0.590 ;
        RECT  6.845 1.310 7.005 1.710 ;
        RECT  6.745 1.550 6.845 1.710 ;
        RECT  6.585 1.550 6.745 2.345 ;
        RECT  5.505 2.185 6.585 2.345 ;
        RECT  6.185 1.685 6.405 1.980 ;
        RECT  6.185 0.770 6.295 0.930 ;
        RECT  6.025 0.770 6.185 1.980 ;
        RECT  5.575 1.165 6.025 1.325 ;
        RECT  5.685 1.505 5.845 2.005 ;
        RECT  5.355 0.770 5.785 0.930 ;
        RECT  5.355 1.505 5.685 1.665 ;
        RECT  5.345 1.845 5.505 2.345 ;
        RECT  5.195 0.770 5.355 1.665 ;
        RECT  2.740 1.845 5.345 2.005 ;
        RECT  4.215 1.505 5.195 1.665 ;
        RECT  4.855 0.430 5.015 1.275 ;
        RECT  4.055 1.015 4.215 1.665 ;
        RECT  4.085 2.185 4.185 2.345 ;
        RECT  3.925 2.185 4.085 2.560 ;
        RECT  3.395 1.505 4.055 1.665 ;
        RECT  2.405 2.400 3.925 2.560 ;
        RECT  3.355 0.345 3.515 0.760 ;
        RECT  3.135 1.320 3.395 1.665 ;
        RECT  1.560 0.345 3.355 0.505 ;
        RECT  2.580 1.785 2.740 2.005 ;
        RECT  1.560 1.785 2.580 1.945 ;
        RECT  2.245 2.125 2.405 2.560 ;
        RECT  0.805 2.125 2.245 2.285 ;
        RECT  1.400 0.345 1.560 1.945 ;
        RECT  1.035 0.720 1.400 0.980 ;
        RECT  1.035 1.685 1.400 1.945 ;
        RECT  0.805 1.175 1.220 1.435 ;
        RECT  0.645 0.680 0.805 2.285 ;
        RECT  0.510 0.680 0.645 0.940 ;
        RECT  0.525 1.795 0.645 2.285 ;
    END
END TLATNSRX1MTH

MACRO TLATNSRX2MTH
    CLASS CORE ;
    FOREIGN TLATNSRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.890 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.150 0.445 1.580 ;
        END
        AntennaGateArea 0.1781 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.925 0.315 6.975 0.475 ;
        RECT  6.765 0.315 6.925 1.305 ;
        RECT  6.715 0.315 6.765 0.475 ;
        RECT  5.335 1.145 6.765 1.305 ;
        RECT  5.175 1.040 5.335 1.305 ;
        RECT  3.730 1.040 5.175 1.200 ;
        RECT  3.570 0.980 3.730 1.200 ;
        RECT  2.915 0.980 3.570 1.140 ;
        RECT  2.815 0.980 2.915 1.170 ;
        RECT  2.655 0.685 2.815 1.170 ;
        RECT  1.950 0.685 2.655 0.845 ;
        RECT  1.790 0.685 1.950 1.580 ;
        RECT  1.740 1.260 1.790 1.580 ;
        END
        AntennaGateArea 0.2535 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.555 0.415 11.790 2.365 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.725 1.290 10.970 1.580 ;
        RECT  10.535 0.765 10.725 2.345 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  9.675 0.880 9.740 1.170 ;
        RECT  9.485 0.880 9.675 1.345 ;
        RECT  9.315 1.185 9.485 1.345 ;
        END
        AntennaGateArea 0.1092 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.435 1.720 4.655 1.880 ;
        RECT  2.150 1.025 2.435 1.880 ;
        END
        AntennaGateArea 0.2834 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.705 -0.130 11.890 0.130 ;
        RECT  9.105 -0.130 9.705 0.250 ;
        RECT  8.665 -0.130 9.105 0.130 ;
        RECT  8.065 -0.130 8.665 0.250 ;
        RECT  6.015 -0.130 8.065 0.130 ;
        RECT  5.855 -0.130 6.015 0.625 ;
        RECT  0.000 -0.130 5.855 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.255 2.740 11.890 3.000 ;
        RECT  10.995 1.845 11.255 3.000 ;
        RECT  9.695 2.740 10.995 3.000 ;
        RECT  9.095 2.480 9.695 3.000 ;
        RECT  7.780 2.740 9.095 3.000 ;
        RECT  7.155 2.245 7.780 3.000 ;
        RECT  5.675 2.740 7.155 3.000 ;
        RECT  5.515 2.525 5.675 3.000 ;
        RECT  0.000 2.740 5.515 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  11.215 0.405 11.375 1.485 ;
        RECT  10.355 0.405 11.215 0.565 ;
        RECT  10.195 0.405 10.355 2.465 ;
        RECT  10.005 0.405 10.195 0.930 ;
        RECT  9.975 1.865 10.195 2.465 ;
        RECT  9.855 1.315 10.015 1.685 ;
        RECT  8.065 0.430 10.005 0.590 ;
        RECT  9.655 1.525 9.855 1.685 ;
        RECT  9.495 1.525 9.655 2.300 ;
        RECT  8.165 2.140 9.495 2.300 ;
        RECT  9.135 0.770 9.305 0.930 ;
        RECT  8.975 0.770 9.135 1.960 ;
        RECT  8.585 1.165 8.975 1.325 ;
        RECT  8.855 1.700 8.975 1.960 ;
        RECT  8.405 0.770 8.795 0.930 ;
        RECT  8.505 1.800 8.605 1.960 ;
        RECT  8.405 1.505 8.505 1.960 ;
        RECT  8.345 0.770 8.405 1.960 ;
        RECT  8.245 0.770 8.345 1.665 ;
        RECT  7.265 1.505 8.245 1.665 ;
        RECT  8.005 1.845 8.165 2.300 ;
        RECT  7.905 0.430 8.065 1.275 ;
        RECT  4.995 1.845 8.005 2.005 ;
        RECT  7.105 1.015 7.265 1.665 ;
        RECT  4.995 1.505 7.105 1.665 ;
        RECT  5.335 2.185 6.745 2.345 ;
        RECT  6.425 0.655 6.585 0.965 ;
        RECT  5.675 0.805 6.425 0.965 ;
        RECT  5.515 0.700 5.675 0.965 ;
        RECT  4.060 0.700 5.515 0.860 ;
        RECT  5.175 2.185 5.335 2.560 ;
        RECT  0.805 2.400 5.175 2.560 ;
        RECT  4.835 1.380 4.995 1.665 ;
        RECT  4.835 1.845 4.995 2.220 ;
        RECT  3.395 1.380 4.835 1.540 ;
        RECT  1.560 2.060 4.835 2.220 ;
        RECT  3.900 0.615 4.060 0.860 ;
        RECT  3.565 0.615 3.900 0.775 ;
        RECT  3.305 0.345 3.565 0.775 ;
        RECT  3.135 1.320 3.395 1.540 ;
        RECT  1.560 0.345 3.305 0.505 ;
        RECT  1.400 0.345 1.560 2.220 ;
        RECT  1.035 0.585 1.400 0.845 ;
        RECT  1.035 1.960 1.400 2.220 ;
        RECT  0.805 1.195 1.220 1.455 ;
        RECT  0.645 0.610 0.805 2.560 ;
        RECT  0.525 0.610 0.645 0.870 ;
        RECT  0.525 1.795 0.645 2.560 ;
    END
END TLATNSRX2MTH

MACRO TLATNSRX4MTH
    CLASS CORE ;
    FOREIGN TLATNSRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.530 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.920 1.235 1.130 1.580 ;
        RECT  0.465 1.235 0.920 1.495 ;
        END
        AntennaGateArea 0.338 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.520 0.315 7.550 0.575 ;
        RECT  7.360 0.315 7.520 1.305 ;
        RECT  5.940 1.145 7.360 1.305 ;
        RECT  5.780 1.040 5.940 1.305 ;
        RECT  4.350 1.040 5.780 1.200 ;
        RECT  4.190 0.980 4.350 1.200 ;
        RECT  3.535 0.980 4.190 1.140 ;
        RECT  3.435 0.980 3.535 1.155 ;
        RECT  3.275 0.685 3.435 1.155 ;
        RECT  2.525 0.685 3.275 0.845 ;
        RECT  2.365 0.685 2.525 1.580 ;
        RECT  2.150 1.150 2.365 1.580 ;
        END
        AntennaGateArea 0.2509 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.965 1.290 13.020 1.580 ;
        RECT  12.765 0.415 12.965 2.365 ;
        RECT  12.650 0.415 12.765 1.015 ;
        RECT  12.635 1.765 12.765 2.365 ;
        END
        AntennaDiffArea 0.684 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.630 0.405 11.890 1.950 ;
        RECT  11.550 1.290 11.630 1.950 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  10.000 0.730 10.245 1.580 ;
        RECT  9.830 1.330 10.000 1.580 ;
        END
        AntennaGateArea 0.1937 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.220 1.720 5.275 1.880 ;
        RECT  3.055 1.330 3.220 1.880 ;
        RECT  2.895 1.025 3.055 1.880 ;
        RECT  2.795 1.025 2.895 1.185 ;
        END
        AntennaGateArea 0.2834 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.400 -0.130 13.530 0.130 ;
        RECT  12.140 -0.130 12.400 1.015 ;
        RECT  11.350 -0.130 12.140 0.130 ;
        RECT  11.090 -0.130 11.350 0.620 ;
        RECT  6.610 -0.130 11.090 0.130 ;
        RECT  6.450 -0.130 6.610 0.625 ;
        RECT  0.385 -0.130 6.450 0.130 ;
        RECT  0.125 -0.130 0.385 0.850 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  13.405 2.740 13.530 3.000 ;
        RECT  13.145 1.845 13.405 3.000 ;
        RECT  10.240 2.740 13.145 3.000 ;
        RECT  9.980 2.545 10.240 3.000 ;
        RECT  8.320 2.740 9.980 3.000 ;
        RECT  7.820 2.245 8.320 3.000 ;
        RECT  6.295 2.740 7.820 3.000 ;
        RECT  6.135 2.525 6.295 3.000 ;
        RECT  0.385 2.740 6.135 3.000 ;
        RECT  0.125 1.755 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.315 1.225 12.585 1.485 ;
        RECT  12.155 1.225 12.315 2.360 ;
        RECT  11.370 2.200 12.155 2.360 ;
        RECT  11.210 0.820 11.370 2.360 ;
        RECT  10.810 0.820 11.210 0.980 ;
        RECT  10.530 2.100 11.210 2.360 ;
        RECT  10.585 1.220 11.025 1.480 ;
        RECT  10.550 0.345 10.810 0.980 ;
        RECT  10.425 1.220 10.585 1.920 ;
        RECT  8.660 0.345 10.550 0.505 ;
        RECT  10.255 1.760 10.425 1.920 ;
        RECT  10.095 1.760 10.255 2.365 ;
        RECT  8.660 2.205 10.095 2.365 ;
        RECT  9.660 0.685 9.820 1.150 ;
        RECT  9.650 1.765 9.705 2.025 ;
        RECT  9.650 0.990 9.660 1.150 ;
        RECT  9.485 0.990 9.650 2.025 ;
        RECT  9.330 1.175 9.485 1.435 ;
        RECT  9.150 0.685 9.310 0.945 ;
        RECT  9.150 1.750 9.190 2.010 ;
        RECT  8.990 0.685 9.150 2.010 ;
        RECT  8.930 1.505 8.990 2.010 ;
        RECT  7.860 1.505 8.930 1.665 ;
        RECT  8.500 0.345 8.660 1.315 ;
        RECT  8.500 1.845 8.660 2.365 ;
        RECT  5.615 1.845 8.500 2.005 ;
        RECT  7.700 1.055 7.860 1.665 ;
        RECT  5.610 1.505 7.700 1.665 ;
        RECT  5.955 2.185 7.340 2.345 ;
        RECT  7.020 0.705 7.180 0.965 ;
        RECT  6.270 0.805 7.020 0.965 ;
        RECT  6.110 0.615 6.270 0.965 ;
        RECT  4.185 0.615 6.110 0.775 ;
        RECT  5.795 2.185 5.955 2.560 ;
        RECT  1.525 2.400 5.795 2.560 ;
        RECT  5.455 1.845 5.615 2.220 ;
        RECT  5.450 1.380 5.610 1.665 ;
        RECT  1.955 2.060 5.455 2.220 ;
        RECT  4.015 1.380 5.450 1.540 ;
        RECT  3.925 0.345 4.185 0.775 ;
        RECT  3.755 1.320 4.015 1.540 ;
        RECT  1.955 0.345 3.925 0.505 ;
        RECT  1.795 0.345 1.955 2.220 ;
        RECT  1.705 0.610 1.795 0.870 ;
        RECT  1.705 1.685 1.795 1.945 ;
        RECT  1.525 1.145 1.615 1.405 ;
        RECT  1.365 0.705 1.525 2.560 ;
        RECT  0.895 0.705 1.365 0.865 ;
        RECT  0.895 2.400 1.365 2.560 ;
        RECT  0.635 0.605 0.895 0.865 ;
        RECT  0.635 1.760 0.895 2.560 ;
    END
END TLATNSRX4MTH

MACRO TLATNTSCAX12MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX12MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.810 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.770 1.115 4.000 1.685 ;
        END
        AntennaGateArea 0.1794 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  16.060 0.485 16.680 2.375 ;
        RECT  12.435 0.485 16.060 0.805 ;
        RECT  15.885 1.400 16.060 2.375 ;
        RECT  15.115 1.905 15.885 2.375 ;
        RECT  12.745 1.905 15.115 2.505 ;
        END
        AntennaDiffArea 1.808 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.095 1.180 3.590 1.580 ;
        END
        AntennaGateArea 0.1794 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.245 1.840 1.540 ;
        END
        AntennaGateArea 0.676 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  16.435 -0.130 16.810 0.130 ;
        RECT  15.835 -0.130 16.435 0.265 ;
        RECT  14.870 -0.130 15.835 0.130 ;
        RECT  14.610 -0.130 14.870 0.265 ;
        RECT  13.645 -0.130 14.610 0.130 ;
        RECT  13.045 -0.130 13.645 0.265 ;
        RECT  10.325 -0.130 13.045 0.130 ;
        RECT  9.725 -0.130 10.325 0.250 ;
        RECT  8.520 -0.130 9.725 0.130 ;
        RECT  7.920 -0.130 8.520 0.250 ;
        RECT  6.975 -0.130 7.920 0.130 ;
        RECT  6.375 -0.130 6.975 0.250 ;
        RECT  3.250 -0.130 6.375 0.130 ;
        RECT  2.990 -0.130 3.250 0.250 ;
        RECT  1.405 -0.130 2.990 0.130 ;
        RECT  1.145 -0.130 1.405 0.720 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.870 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  15.610 2.740 16.810 3.000 ;
        RECT  15.350 2.595 15.610 3.000 ;
        RECT  12.085 2.740 15.350 3.000 ;
        RECT  11.585 2.195 12.085 3.000 ;
        RECT  8.525 2.740 11.585 3.000 ;
        RECT  7.925 2.620 8.525 3.000 ;
        RECT  6.975 2.740 7.925 3.000 ;
        RECT  6.375 2.620 6.975 3.000 ;
        RECT  5.285 2.740 6.375 3.000 ;
        RECT  5.025 2.620 5.285 3.000 ;
        RECT  2.335 2.740 5.025 3.000 ;
        RECT  2.075 2.105 2.335 3.000 ;
        RECT  0.385 2.740 2.075 3.000 ;
        RECT  0.125 1.720 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  15.675 1.055 15.880 1.215 ;
        RECT  15.515 1.055 15.675 1.685 ;
        RECT  14.855 1.525 15.515 1.685 ;
        RECT  15.075 1.025 15.335 1.345 ;
        RECT  13.995 1.025 15.075 1.185 ;
        RECT  14.255 1.365 14.855 1.685 ;
        RECT  13.175 1.525 14.255 1.685 ;
        RECT  13.395 1.025 13.995 1.345 ;
        RECT  12.300 1.025 13.395 1.185 ;
        RECT  12.575 1.365 13.175 1.685 ;
        RECT  11.860 1.525 12.575 1.685 ;
        RECT  12.200 1.025 12.300 1.345 ;
        RECT  12.040 0.310 12.200 1.345 ;
        RECT  10.695 0.310 12.040 0.470 ;
        RECT  11.700 0.650 11.860 1.945 ;
        RECT  11.030 0.650 11.700 0.810 ;
        RECT  11.560 1.685 11.700 1.945 ;
        RECT  11.370 1.005 11.520 1.265 ;
        RECT  11.210 1.005 11.370 2.560 ;
        RECT  9.300 2.400 11.210 2.560 ;
        RECT  10.870 0.650 11.030 2.220 ;
        RECT  10.070 2.060 10.870 2.220 ;
        RECT  10.535 0.310 10.695 0.590 ;
        RECT  10.505 0.775 10.690 1.860 ;
        RECT  9.300 0.430 10.535 0.590 ;
        RECT  10.250 0.775 10.505 0.935 ;
        RECT  10.250 1.700 10.505 1.860 ;
        RECT  10.070 1.205 10.210 1.465 ;
        RECT  9.910 0.810 10.070 2.220 ;
        RECT  5.770 0.810 9.910 0.970 ;
        RECT  5.770 1.755 9.910 1.915 ;
        RECT  9.570 1.205 9.730 1.465 ;
        RECT  5.330 1.285 9.570 1.465 ;
        RECT  8.700 0.310 9.300 0.590 ;
        RECT  8.700 2.100 9.300 2.560 ;
        RECT  7.750 0.430 8.700 0.590 ;
        RECT  7.750 2.100 8.700 2.260 ;
        RECT  7.150 0.310 7.750 0.590 ;
        RECT  7.150 2.100 7.750 2.560 ;
        RECT  6.200 0.430 7.150 0.590 ;
        RECT  6.200 2.100 7.150 2.260 ;
        RECT  5.760 0.310 6.200 0.590 ;
        RECT  5.600 2.100 6.200 2.560 ;
        RECT  5.600 0.310 5.760 0.565 ;
        RECT  4.345 0.405 5.600 0.565 ;
        RECT  2.865 2.210 5.600 2.370 ;
        RECT  5.170 0.865 5.330 2.005 ;
        RECT  4.680 0.865 5.170 1.025 ;
        RECT  4.680 1.845 5.170 2.005 ;
        RECT  4.340 1.210 4.900 1.470 ;
        RECT  4.520 0.765 4.680 1.025 ;
        RECT  4.520 1.685 4.680 2.005 ;
        RECT  4.185 0.405 4.345 0.590 ;
        RECT  4.180 0.775 4.340 2.030 ;
        RECT  2.400 0.430 4.185 0.590 ;
        RECT  3.530 0.775 4.180 0.935 ;
        RECT  3.095 1.870 4.180 2.030 ;
        RECT  2.705 0.815 2.865 2.370 ;
        RECT  2.595 0.815 2.705 0.975 ;
        RECT  2.585 1.770 2.705 2.370 ;
        RECT  2.400 1.245 2.515 1.505 ;
        RECT  2.240 0.430 2.400 1.880 ;
        RECT  1.915 0.900 2.240 1.060 ;
        RECT  1.825 1.720 2.240 1.880 ;
        RECT  1.655 0.655 1.915 1.060 ;
        RECT  1.565 1.720 1.825 2.325 ;
        RECT  0.895 0.900 1.655 1.060 ;
        RECT  0.895 1.720 1.565 1.880 ;
        RECT  0.635 0.660 0.895 1.060 ;
        RECT  0.635 1.720 0.895 2.330 ;
    END
END TLATNTSCAX12MTH

MACRO TLATNTSCAX16MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX16MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 22.550 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.575 1.250 4.000 1.635 ;
        END
        AntennaGateArea 0.2366 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  19.825 0.810 22.425 1.100 ;
        RECT  19.825 1.660 22.090 2.060 ;
        RECT  19.125 0.810 19.825 2.060 ;
        RECT  16.220 0.810 19.125 1.100 ;
        RECT  16.640 1.660 19.125 2.060 ;
        END
        AntennaDiffArea 2.862 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.180 1.180 4.770 1.630 ;
        END
        AntennaGateArea 0.2366 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.505 1.290 2.465 1.540 ;
        END
        AntennaGateArea 0.8658 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.885 -0.130 22.550 0.130 ;
        RECT  21.625 -0.130 21.885 0.590 ;
        RECT  20.250 -0.130 21.625 0.130 ;
        RECT  19.990 -0.130 20.250 0.250 ;
        RECT  18.695 -0.130 19.990 0.130 ;
        RECT  17.755 -0.130 18.695 0.250 ;
        RECT  17.020 -0.130 17.755 0.130 ;
        RECT  16.760 -0.130 17.020 0.250 ;
        RECT  14.110 -0.130 16.760 0.130 ;
        RECT  13.510 -0.130 14.110 0.250 ;
        RECT  12.070 -0.130 13.510 0.130 ;
        RECT  11.810 -0.130 12.070 0.250 ;
        RECT  10.670 -0.130 11.810 0.130 ;
        RECT  10.410 -0.130 10.670 0.250 ;
        RECT  9.110 -0.130 10.410 0.130 ;
        RECT  8.850 -0.130 9.110 0.250 ;
        RECT  7.550 -0.130 8.850 0.130 ;
        RECT  7.290 -0.130 7.550 0.250 ;
        RECT  5.560 -0.130 7.290 0.130 ;
        RECT  4.960 -0.130 5.560 0.250 ;
        RECT  4.450 -0.130 4.960 0.130 ;
        RECT  3.850 -0.130 4.450 0.250 ;
        RECT  3.615 -0.130 3.850 0.130 ;
        RECT  2.675 -0.130 3.615 0.250 ;
        RECT  0.895 -0.130 2.675 0.130 ;
        RECT  0.635 -0.130 0.895 0.680 ;
        RECT  0.000 -0.130 0.635 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  21.290 2.740 22.550 3.000 ;
        RECT  21.030 2.620 21.290 3.000 ;
        RECT  19.575 2.740 21.030 3.000 ;
        RECT  19.315 2.620 19.575 3.000 ;
        RECT  17.785 2.740 19.315 3.000 ;
        RECT  17.525 2.620 17.785 3.000 ;
        RECT  16.050 2.740 17.525 3.000 ;
        RECT  15.450 2.620 16.050 3.000 ;
        RECT  12.315 2.740 15.450 3.000 ;
        RECT  11.715 2.620 12.315 3.000 ;
        RECT  10.760 2.740 11.715 3.000 ;
        RECT  10.160 2.620 10.760 3.000 ;
        RECT  9.200 2.740 10.160 3.000 ;
        RECT  8.600 2.620 9.200 3.000 ;
        RECT  7.410 2.740 8.600 3.000 ;
        RECT  7.150 2.620 7.410 3.000 ;
        RECT  5.500 2.740 7.150 3.000 ;
        RECT  5.240 2.620 5.500 3.000 ;
        RECT  3.635 2.740 5.240 3.000 ;
        RECT  2.675 2.600 3.635 3.000 ;
        RECT  0.895 2.740 2.675 3.000 ;
        RECT  0.635 2.105 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  22.270 1.280 22.430 2.440 ;
        RECT  20.225 1.280 22.270 1.440 ;
        RECT  16.460 2.280 22.270 2.440 ;
        RECT  20.825 0.310 21.085 0.590 ;
        RECT  19.410 0.430 20.825 0.590 ;
        RECT  19.150 0.310 19.410 0.590 ;
        RECT  17.580 0.430 19.150 0.590 ;
        RECT  16.460 1.280 18.850 1.440 ;
        RECT  17.320 0.310 17.580 0.590 ;
        RECT  16.040 0.430 17.320 0.590 ;
        RECT  16.300 1.280 16.460 2.440 ;
        RECT  15.700 2.280 16.300 2.440 ;
        RECT  15.880 0.310 16.040 1.505 ;
        RECT  14.450 0.310 15.880 0.470 ;
        RECT  15.540 0.650 15.700 2.440 ;
        RECT  14.820 0.650 15.540 0.810 ;
        RECT  15.350 1.685 15.540 1.945 ;
        RECT  15.160 1.020 15.360 1.180 ;
        RECT  15.000 1.020 15.160 2.560 ;
        RECT  13.090 2.400 15.000 2.560 ;
        RECT  14.660 0.650 14.820 2.220 ;
        RECT  13.860 2.060 14.660 2.220 ;
        RECT  14.340 1.245 14.480 1.505 ;
        RECT  14.290 0.310 14.450 0.590 ;
        RECT  14.180 0.775 14.340 1.860 ;
        RECT  13.090 0.430 14.290 0.590 ;
        RECT  14.040 0.775 14.180 0.935 ;
        RECT  14.040 1.700 14.180 1.860 ;
        RECT  13.860 1.205 14.000 1.465 ;
        RECT  13.700 0.810 13.860 2.220 ;
        RECT  8.000 0.810 13.700 0.970 ;
        RECT  8.000 1.755 13.700 1.915 ;
        RECT  13.360 1.205 13.520 1.465 ;
        RECT  7.040 1.285 13.360 1.465 ;
        RECT  12.490 0.310 13.090 0.590 ;
        RECT  12.490 2.100 13.090 2.560 ;
        RECT  11.540 0.430 12.490 0.590 ;
        RECT  11.540 2.100 12.490 2.260 ;
        RECT  10.940 0.310 11.540 0.590 ;
        RECT  10.940 2.100 11.540 2.560 ;
        RECT  9.990 0.430 10.940 0.590 ;
        RECT  9.990 2.100 10.940 2.260 ;
        RECT  9.390 0.310 9.990 0.590 ;
        RECT  9.390 2.100 9.990 2.560 ;
        RECT  8.430 0.430 9.390 0.590 ;
        RECT  8.430 2.100 9.390 2.260 ;
        RECT  7.830 0.310 8.430 0.590 ;
        RECT  7.830 2.100 8.430 2.560 ;
        RECT  2.805 0.430 7.830 0.590 ;
        RECT  3.395 2.210 7.830 2.370 ;
        RECT  6.880 0.815 7.040 2.005 ;
        RECT  5.840 0.815 6.880 0.975 ;
        RECT  5.760 1.845 6.880 2.005 ;
        RECT  5.160 1.210 6.620 1.470 ;
        RECT  5.000 0.815 5.160 2.030 ;
        RECT  3.955 0.815 5.000 0.975 ;
        RECT  4.360 1.870 5.000 2.030 ;
        RECT  3.235 0.815 3.395 2.370 ;
        RECT  3.015 0.815 3.235 0.975 ;
        RECT  3.015 1.805 3.235 2.065 ;
        RECT  2.805 1.245 3.055 1.505 ;
        RECT  2.645 0.430 2.805 1.920 ;
        RECT  2.335 0.865 2.645 1.025 ;
        RECT  2.335 1.760 2.645 1.920 ;
        RECT  2.075 0.605 2.335 1.025 ;
        RECT  2.075 1.760 2.335 2.345 ;
        RECT  1.405 0.865 2.075 1.025 ;
        RECT  1.405 1.760 2.075 1.920 ;
        RECT  1.145 0.605 1.405 1.025 ;
        RECT  1.145 1.760 1.405 2.360 ;
        RECT  0.385 0.865 1.145 1.025 ;
        RECT  0.385 1.760 1.145 1.920 ;
        RECT  0.125 0.605 0.385 1.025 ;
        RECT  0.125 1.760 0.385 2.360 ;
    END
END TLATNTSCAX16MTH

MACRO TLATNTSCAX20MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX20MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 25.010 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.760 1.205 4.195 1.725 ;
        END
        AntennaGateArea 0.2574 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  23.825 0.480 24.665 2.395 ;
        RECT  16.955 0.480 23.825 0.770 ;
        RECT  23.415 1.490 23.825 2.395 ;
        RECT  16.535 2.015 23.415 2.395 ;
        END
        AntennaDiffArea 2.79 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.375 1.180 4.820 1.630 ;
        END
        AntennaGateArea 0.2574 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.550 1.290 2.510 1.540 ;
        END
        AntennaGateArea 1.027 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.595 -0.130 25.010 0.130 ;
        RECT  24.335 -0.130 24.595 0.300 ;
        RECT  23.995 -0.130 24.335 0.130 ;
        RECT  23.055 -0.130 23.995 0.300 ;
        RECT  22.175 -0.130 23.055 0.130 ;
        RECT  21.575 -0.130 22.175 0.300 ;
        RECT  20.635 -0.130 21.575 0.130 ;
        RECT  20.035 -0.130 20.635 0.300 ;
        RECT  19.175 -0.130 20.035 0.130 ;
        RECT  18.575 -0.130 19.175 0.300 ;
        RECT  17.755 -0.130 18.575 0.130 ;
        RECT  17.495 -0.130 17.755 0.300 ;
        RECT  16.675 -0.130 17.495 0.130 ;
        RECT  16.415 -0.130 16.675 0.295 ;
        RECT  12.630 -0.130 16.415 0.130 ;
        RECT  12.370 -0.130 12.630 0.250 ;
        RECT  11.505 -0.130 12.370 0.130 ;
        RECT  11.245 -0.130 11.505 0.250 ;
        RECT  9.950 -0.130 11.245 0.130 ;
        RECT  9.690 -0.130 9.950 0.250 ;
        RECT  8.530 -0.130 9.690 0.130 ;
        RECT  8.270 -0.130 8.530 0.250 ;
        RECT  5.690 -0.130 8.270 0.130 ;
        RECT  5.090 -0.130 5.690 0.295 ;
        RECT  4.820 -0.130 5.090 0.130 ;
        RECT  4.560 -0.130 4.820 0.295 ;
        RECT  4.300 -0.130 4.560 0.130 ;
        RECT  3.700 -0.130 4.300 0.295 ;
        RECT  2.880 -0.130 3.700 0.130 ;
        RECT  2.620 -0.130 2.880 0.295 ;
        RECT  0.900 -0.130 2.620 0.130 ;
        RECT  0.640 -0.130 0.900 0.685 ;
        RECT  0.000 -0.130 0.640 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  24.475 2.740 25.010 3.000 ;
        RECT  23.875 2.620 24.475 3.000 ;
        RECT  20.875 2.740 23.875 3.000 ;
        RECT  20.615 2.575 20.875 3.000 ;
        RECT  17.605 2.740 20.615 3.000 ;
        RECT  17.345 2.575 17.605 3.000 ;
        RECT  15.665 2.740 17.345 3.000 ;
        RECT  15.405 2.610 15.665 3.000 ;
        RECT  14.735 2.740 15.405 3.000 ;
        RECT  14.515 2.100 14.735 3.000 ;
        RECT  13.250 2.740 14.515 3.000 ;
        RECT  12.650 2.620 13.250 3.000 ;
        RECT  11.530 2.740 12.650 3.000 ;
        RECT  11.270 2.620 11.530 3.000 ;
        RECT  9.980 2.740 11.270 3.000 ;
        RECT  9.720 2.620 9.980 3.000 ;
        RECT  8.420 2.740 9.720 3.000 ;
        RECT  8.160 2.620 8.420 3.000 ;
        RECT  3.845 2.740 8.160 3.000 ;
        RECT  3.585 2.580 3.845 3.000 ;
        RECT  2.880 2.740 3.585 3.000 ;
        RECT  2.620 2.555 2.880 3.000 ;
        RECT  0.900 2.740 2.620 3.000 ;
        RECT  0.640 2.105 0.900 3.000 ;
        RECT  0.000 2.740 0.640 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  23.375 0.955 23.605 1.215 ;
        RECT  22.565 0.955 23.375 1.115 ;
        RECT  22.855 1.320 23.115 1.795 ;
        RECT  21.895 1.635 22.855 1.795 ;
        RECT  22.305 0.955 22.565 1.455 ;
        RECT  21.035 0.955 22.305 1.115 ;
        RECT  21.295 1.295 21.895 1.795 ;
        RECT  20.195 1.635 21.295 1.795 ;
        RECT  20.435 0.955 21.035 1.455 ;
        RECT  19.300 0.955 20.435 1.115 ;
        RECT  19.595 1.295 20.195 1.795 ;
        RECT  18.635 1.635 19.595 1.795 ;
        RECT  19.040 0.955 19.300 1.455 ;
        RECT  17.765 0.955 19.040 1.115 ;
        RECT  18.300 1.295 18.635 1.795 ;
        RECT  16.915 1.635 18.300 1.795 ;
        RECT  17.165 0.955 17.765 1.420 ;
        RECT  16.585 0.955 17.165 1.115 ;
        RECT  16.655 1.315 16.915 1.795 ;
        RECT  16.425 0.475 16.585 1.115 ;
        RECT  16.235 0.475 16.425 0.635 ;
        RECT  16.245 1.325 16.325 2.430 ;
        RECT  16.165 0.815 16.245 2.430 ;
        RECT  16.075 0.310 16.235 0.635 ;
        RECT  16.085 0.815 16.165 1.485 ;
        RECT  15.175 2.270 16.165 2.430 ;
        RECT  15.985 0.815 16.085 0.975 ;
        RECT  12.970 0.310 16.075 0.470 ;
        RECT  15.825 1.760 15.985 2.070 ;
        RECT  15.805 1.760 15.825 1.920 ;
        RECT  15.645 0.700 15.805 1.920 ;
        RECT  13.310 0.700 15.645 0.860 ;
        RECT  13.920 1.760 15.645 1.920 ;
        RECT  15.365 1.070 15.465 1.230 ;
        RECT  15.205 1.070 15.365 1.545 ;
        RECT  13.830 1.385 15.205 1.545 ;
        RECT  14.915 2.270 15.175 2.510 ;
        RECT  13.650 1.045 14.665 1.205 ;
        RECT  13.490 2.280 14.090 2.560 ;
        RECT  13.660 1.760 13.920 2.095 ;
        RECT  12.230 1.760 13.660 1.920 ;
        RECT  13.490 1.045 13.650 1.455 ;
        RECT  7.050 1.295 13.490 1.455 ;
        RECT  12.400 2.280 13.490 2.440 ;
        RECT  13.150 0.700 13.310 1.075 ;
        RECT  12.365 0.915 13.150 1.075 ;
        RECT  12.810 0.310 12.970 0.640 ;
        RECT  12.190 0.480 12.810 0.640 ;
        RECT  11.800 2.280 12.400 2.560 ;
        RECT  12.105 0.820 12.365 1.075 ;
        RECT  11.970 1.760 12.230 2.095 ;
        RECT  11.935 0.310 12.190 0.640 ;
        RECT  10.800 0.915 12.105 1.075 ;
        RECT  10.680 1.760 11.970 1.920 ;
        RECT  11.930 0.310 11.935 0.590 ;
        RECT  10.970 0.430 11.930 0.590 ;
        RECT  10.850 2.280 11.800 2.440 ;
        RECT  10.370 0.310 10.970 0.590 ;
        RECT  10.250 2.280 10.850 2.560 ;
        RECT  10.540 0.770 10.800 1.075 ;
        RECT  10.420 1.760 10.680 2.095 ;
        RECT  9.240 0.915 10.540 1.075 ;
        RECT  9.130 1.760 10.420 1.920 ;
        RECT  9.410 0.430 10.370 0.590 ;
        RECT  9.300 2.280 10.250 2.440 ;
        RECT  8.810 0.310 9.410 0.590 ;
        RECT  8.700 2.280 9.300 2.560 ;
        RECT  8.980 0.770 9.240 1.075 ;
        RECT  8.870 1.760 9.130 2.095 ;
        RECT  7.680 0.915 8.980 1.075 ;
        RECT  7.570 1.760 8.870 1.920 ;
        RECT  7.420 0.430 8.810 0.590 ;
        RECT  7.310 2.280 8.700 2.440 ;
        RECT  7.420 0.770 7.680 1.075 ;
        RECT  7.310 1.760 7.570 2.060 ;
        RECT  7.160 0.310 7.420 0.590 ;
        RECT  7.050 2.240 7.310 2.560 ;
        RECT  6.055 0.430 7.160 0.590 ;
        RECT  7.050 0.815 7.160 0.975 ;
        RECT  6.890 0.815 7.050 2.060 ;
        RECT  3.580 2.240 7.050 2.400 ;
        RECT  5.970 0.815 6.890 0.975 ;
        RECT  6.790 1.800 6.890 2.060 ;
        RECT  6.110 1.800 6.790 1.960 ;
        RECT  5.290 1.265 6.710 1.425 ;
        RECT  5.850 1.800 6.110 2.060 ;
        RECT  5.895 0.430 6.055 0.635 ;
        RECT  2.895 0.475 5.895 0.635 ;
        RECT  5.130 0.815 5.290 2.030 ;
        RECT  4.100 0.815 5.130 0.975 ;
        RECT  4.460 1.870 5.130 2.030 ;
        RECT  3.420 0.815 3.580 2.400 ;
        RECT  3.160 0.815 3.420 0.975 ;
        RECT  3.075 1.830 3.420 2.090 ;
        RECT  2.895 1.245 3.240 1.505 ;
        RECT  2.735 0.475 2.895 1.920 ;
        RECT  2.340 0.865 2.735 1.025 ;
        RECT  2.340 1.760 2.735 1.920 ;
        RECT  2.080 0.425 2.340 1.025 ;
        RECT  2.080 1.760 2.340 2.415 ;
        RECT  1.410 0.865 2.080 1.025 ;
        RECT  1.410 1.760 2.080 1.920 ;
        RECT  1.150 0.425 1.410 1.025 ;
        RECT  1.150 1.760 1.410 2.415 ;
        RECT  0.390 0.865 1.150 1.025 ;
        RECT  0.390 1.760 1.150 1.920 ;
        RECT  0.130 0.425 0.390 1.025 ;
        RECT  0.130 1.760 0.390 2.415 ;
    END
END TLATNTSCAX20MTH

MACRO TLATNTSCAX2MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.970 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.270 0.450 1.715 ;
        END
        AntennaGateArea 0.0624 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.660 0.815 6.870 2.415 ;
        RECT  6.045 0.815 6.660 0.975 ;
        RECT  6.585 1.815 6.660 2.415 ;
        END
        AntennaDiffArea 0.414 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.455 2.075 0.905 2.380 ;
        END
        AntennaGateArea 0.0624 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  1.740 1.350 2.015 1.990 ;
        END
        AntennaGateArea 0.1391 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.845 -0.130 6.970 0.130 ;
        RECT  6.585 -0.130 6.845 0.635 ;
        RECT  6.005 -0.130 6.585 0.130 ;
        RECT  5.065 -0.130 6.005 0.250 ;
        RECT  3.435 -0.130 5.065 0.130 ;
        RECT  3.175 -0.130 3.435 0.605 ;
        RECT  1.385 -0.130 3.175 0.130 ;
        RECT  1.125 -0.130 1.385 0.505 ;
        RECT  0.385 -0.130 1.125 0.130 ;
        RECT  0.125 -0.130 0.385 0.380 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.895 2.740 6.970 3.000 ;
        RECT  5.295 2.540 5.895 3.000 ;
        RECT  3.360 2.740 5.295 3.000 ;
        RECT  2.760 2.510 3.360 3.000 ;
        RECT  1.835 2.740 2.760 3.000 ;
        RECT  1.575 2.410 1.835 3.000 ;
        RECT  0.385 2.740 1.575 3.000 ;
        RECT  0.125 2.560 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.235 0.330 6.395 0.590 ;
        RECT  4.855 0.430 6.235 0.590 ;
        RECT  6.070 1.300 6.115 1.560 ;
        RECT  5.910 1.300 6.070 2.360 ;
        RECT  4.735 2.200 5.910 2.360 ;
        RECT  5.570 0.815 5.730 1.915 ;
        RECT  5.065 0.815 5.570 0.975 ;
        RECT  4.825 1.735 5.570 1.915 ;
        RECT  4.395 1.275 5.390 1.435 ;
        RECT  4.695 0.430 4.855 0.895 ;
        RECT  4.575 2.200 4.735 2.560 ;
        RECT  4.395 0.735 4.695 0.895 ;
        RECT  3.710 2.400 4.575 2.560 ;
        RECT  3.775 0.310 4.515 0.470 ;
        RECT  4.235 0.735 4.395 2.190 ;
        RECT  3.995 0.735 4.235 0.895 ;
        RECT  3.950 1.930 4.235 2.190 ;
        RECT  3.895 1.080 4.055 1.340 ;
        RECT  3.440 1.180 3.895 1.340 ;
        RECT  3.615 0.310 3.775 0.945 ;
        RECT  3.550 2.170 3.710 2.560 ;
        RECT  2.865 0.785 3.615 0.945 ;
        RECT  3.440 2.170 3.550 2.330 ;
        RECT  3.280 1.180 3.440 2.330 ;
        RECT  2.375 2.170 3.280 2.330 ;
        RECT  2.705 0.785 2.865 1.990 ;
        RECT  1.725 0.310 2.790 0.470 ;
        RECT  2.605 0.785 2.705 0.975 ;
        RECT  2.565 1.730 2.705 1.990 ;
        RECT  2.355 1.300 2.505 1.560 ;
        RECT  2.355 2.170 2.375 2.515 ;
        RECT  2.195 0.765 2.355 2.515 ;
        RECT  2.145 0.765 2.195 1.025 ;
        RECT  2.115 2.170 2.195 2.515 ;
        RECT  1.565 0.310 1.725 0.925 ;
        RECT  1.525 0.765 1.565 0.925 ;
        RECT  1.365 0.765 1.525 2.235 ;
        RECT  1.125 0.765 1.365 1.025 ;
        RECT  1.245 2.075 1.365 2.235 ;
        RECT  1.085 2.075 1.245 2.515 ;
        RECT  0.880 1.265 1.185 1.525 ;
        RECT  0.880 1.735 1.095 1.895 ;
        RECT  0.720 0.585 0.880 1.895 ;
        RECT  0.555 0.585 0.720 0.845 ;
    END
END TLATNTSCAX2MTH

MACRO TLATNTSCAX3MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.325 1.025 0.585 1.580 ;
        RECT  0.100 1.290 0.325 1.580 ;
        END
        AntennaGateArea 0.0624 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.400 0.555 7.530 0.815 ;
        RECT  7.150 0.555 7.400 1.990 ;
        RECT  6.930 1.700 7.150 1.990 ;
        END
        AntennaDiffArea 0.428 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.645 2.095 1.220 2.400 ;
        END
        AntennaGateArea 0.0624 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  2.085 1.305 2.390 1.990 ;
        END
        AntennaGateArea 0.1846 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.075 -0.130 8.200 0.130 ;
        RECT  7.815 -0.130 8.075 0.825 ;
        RECT  5.660 -0.130 7.815 0.130 ;
        RECT  5.460 -0.130 5.660 0.435 ;
        RECT  4.080 -0.130 5.460 0.130 ;
        RECT  3.820 -0.130 4.080 0.250 ;
        RECT  2.010 -0.130 3.820 0.130 ;
        RECT  1.410 -0.130 2.010 0.425 ;
        RECT  0.385 -0.130 1.410 0.130 ;
        RECT  0.125 -0.130 0.385 0.845 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.060 2.740 8.200 3.000 ;
        RECT  7.800 2.550 8.060 3.000 ;
        RECT  6.220 2.740 7.800 3.000 ;
        RECT  5.280 2.550 6.220 3.000 ;
        RECT  3.750 2.740 5.280 3.000 ;
        RECT  3.150 2.550 3.750 3.000 ;
        RECT  2.285 2.740 3.150 3.000 ;
        RECT  2.025 2.230 2.285 3.000 ;
        RECT  1.660 2.740 2.025 3.000 ;
        RECT  0.720 2.620 1.660 3.000 ;
        RECT  0.385 2.740 0.720 3.000 ;
        RECT  0.125 1.940 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.740 1.155 7.840 1.415 ;
        RECT  7.580 1.155 7.740 2.350 ;
        RECT  6.490 2.190 7.580 2.350 ;
        RECT  6.810 0.310 6.970 1.380 ;
        RECT  6.010 0.310 6.810 0.470 ;
        RECT  6.330 1.315 6.490 2.350 ;
        RECT  6.190 0.685 6.450 1.135 ;
        RECT  4.970 2.190 6.330 2.350 ;
        RECT  6.115 0.975 6.190 1.135 ;
        RECT  5.955 0.975 6.115 1.470 ;
        RECT  5.850 0.310 6.010 0.775 ;
        RECT  5.860 1.310 5.955 1.470 ;
        RECT  5.600 1.310 5.860 1.945 ;
        RECT  5.685 0.615 5.850 0.775 ;
        RECT  5.525 0.615 5.685 0.845 ;
        RECT  5.410 1.310 5.600 1.570 ;
        RECT  4.830 0.685 5.525 0.845 ;
        RECT  4.420 0.310 5.190 0.470 ;
        RECT  4.710 2.190 4.970 2.485 ;
        RECT  4.670 0.685 4.830 1.915 ;
        RECT  2.900 2.190 4.710 2.350 ;
        RECT  4.340 1.755 4.670 1.915 ;
        RECT  4.260 0.310 4.420 1.575 ;
        RECT  3.510 0.430 4.260 0.590 ;
        RECT  4.160 1.315 4.260 1.575 ;
        RECT  4.000 1.315 4.160 1.865 ;
        RECT  3.240 1.705 4.000 1.865 ;
        RECT  3.660 0.855 3.820 1.265 ;
        RECT  3.070 0.855 3.660 1.015 ;
        RECT  3.250 0.360 3.510 0.590 ;
        RECT  2.900 1.200 3.390 1.460 ;
        RECT  3.080 1.705 3.240 1.965 ;
        RECT  2.910 0.425 3.070 1.015 ;
        RECT  2.385 0.425 2.910 0.585 ;
        RECT  2.740 1.200 2.900 2.425 ;
        RECT  2.730 1.200 2.740 1.460 ;
        RECT  2.580 2.165 2.740 2.425 ;
        RECT  2.570 0.765 2.730 1.460 ;
        RECT  2.225 0.425 2.385 0.925 ;
        RECT  1.760 0.765 2.225 0.925 ;
        RECT  1.600 0.765 1.760 2.010 ;
        RECT  1.485 0.765 1.600 1.025 ;
        RECT  1.485 1.750 1.600 2.010 ;
        RECT  0.995 1.265 1.405 1.525 ;
        RECT  0.995 1.735 1.235 1.895 ;
        RECT  0.835 0.480 0.995 1.895 ;
        RECT  0.695 0.480 0.835 0.740 ;
    END
END TLATNTSCAX3MTH

MACRO TLATNTSCAX4MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.155 2.975 1.580 ;
        END
        AntennaGateArea 0.0806 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.560 0.600 9.740 2.045 ;
        RECT  8.525 0.600 9.560 0.780 ;
        RECT  9.445 1.600 9.560 2.045 ;
        RECT  8.835 1.865 9.445 2.045 ;
        RECT  8.575 1.865 8.835 2.465 ;
        RECT  8.265 0.520 8.525 0.780 ;
        END
        AntennaDiffArea 0.572 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 1.095 2.380 1.580 ;
        END
        AntennaGateArea 0.0806 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 1.035 1.465 ;
        RECT  0.100 1.205 0.310 1.705 ;
        END
        AntennaGateArea 0.2392 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.455 -0.130 9.840 0.130 ;
        RECT  8.855 -0.130 9.455 0.315 ;
        RECT  6.160 -0.130 8.855 0.130 ;
        RECT  5.560 -0.130 6.160 0.250 ;
        RECT  2.705 -0.130 5.560 0.130 ;
        RECT  1.765 -0.130 2.705 0.250 ;
        RECT  1.545 -0.130 1.765 0.130 ;
        RECT  0.605 -0.130 1.545 0.250 ;
        RECT  0.425 -0.130 0.605 0.130 ;
        RECT  0.165 -0.130 0.425 0.970 ;
        RECT  0.000 -0.130 0.165 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.655 2.740 9.840 3.000 ;
        RECT  9.395 2.225 9.655 3.000 ;
        RECT  7.925 2.740 9.395 3.000 ;
        RECT  7.425 2.195 7.925 3.000 ;
        RECT  4.110 2.740 7.425 3.000 ;
        RECT  3.170 2.620 4.110 3.000 ;
        RECT  2.740 2.740 3.170 3.000 ;
        RECT  1.800 2.620 2.740 3.000 ;
        RECT  1.325 2.740 1.800 3.000 ;
        RECT  1.065 1.985 1.325 3.000 ;
        RECT  0.770 2.740 1.065 3.000 ;
        RECT  0.170 2.480 0.770 3.000 ;
        RECT  0.000 2.740 0.170 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.055 1.000 9.315 1.260 ;
        RECT  8.185 1.000 9.055 1.160 ;
        RECT  8.405 1.365 8.665 1.685 ;
        RECT  7.700 1.525 8.405 1.685 ;
        RECT  8.080 1.000 8.185 1.325 ;
        RECT  7.920 0.310 8.080 1.325 ;
        RECT  6.535 0.310 7.920 0.470 ;
        RECT  7.540 0.650 7.700 1.945 ;
        RECT  6.870 0.650 7.540 0.810 ;
        RECT  7.400 1.685 7.540 1.945 ;
        RECT  7.210 1.005 7.360 1.265 ;
        RECT  7.050 1.005 7.210 2.560 ;
        RECT  5.140 2.400 7.050 2.560 ;
        RECT  6.710 0.650 6.870 2.220 ;
        RECT  5.910 2.060 6.710 2.220 ;
        RECT  6.375 0.310 6.535 0.590 ;
        RECT  6.345 0.785 6.530 1.865 ;
        RECT  5.140 0.430 6.375 0.590 ;
        RECT  6.090 0.785 6.345 0.945 ;
        RECT  6.090 1.705 6.345 1.865 ;
        RECT  5.910 1.215 6.050 1.475 ;
        RECT  5.750 0.810 5.910 2.220 ;
        RECT  4.710 0.810 5.750 0.970 ;
        RECT  4.970 1.800 5.750 1.960 ;
        RECT  3.845 1.235 5.570 1.495 ;
        RECT  4.540 0.310 5.140 0.590 ;
        RECT  4.540 2.280 5.140 2.560 ;
        RECT  4.710 1.800 4.970 2.060 ;
        RECT  4.140 0.430 4.540 0.590 ;
        RECT  1.885 2.280 4.540 2.440 ;
        RECT  3.980 0.405 4.140 0.590 ;
        RECT  3.365 0.405 3.980 0.565 ;
        RECT  3.685 0.765 3.845 1.950 ;
        RECT  3.540 0.765 3.685 1.025 ;
        RECT  3.540 1.690 3.685 1.950 ;
        RECT  3.360 1.235 3.505 1.495 ;
        RECT  3.205 0.405 3.365 0.590 ;
        RECT  3.200 0.815 3.360 1.920 ;
        RECT  1.420 0.430 3.205 0.590 ;
        RECT  2.550 0.815 3.200 0.975 ;
        RECT  2.115 1.760 3.200 1.920 ;
        RECT  1.725 0.815 1.885 2.440 ;
        RECT  1.615 0.815 1.725 0.975 ;
        RECT  1.605 1.685 1.725 2.440 ;
        RECT  1.420 1.205 1.545 1.465 ;
        RECT  1.260 0.430 1.420 1.805 ;
        RECT  0.675 0.710 1.260 0.970 ;
        RECT  0.785 1.645 1.260 1.805 ;
        RECT  0.525 1.645 0.785 2.060 ;
    END
END TLATNTSCAX4MTH

MACRO TLATNTSCAX6MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX6MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.155 2.975 1.635 ;
        END
        AntennaGateArea 0.0988 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  11.110 0.555 11.380 2.465 ;
        RECT  9.110 0.555 11.110 0.825 ;
        RECT  11.095 1.855 11.110 2.465 ;
        RECT  9.675 1.855 11.095 2.125 ;
        RECT  9.415 1.855 9.675 2.465 ;
        END
        AntennaDiffArea 1.018 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 1.120 2.380 1.680 ;
        END
        AntennaGateArea 0.0988 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 0.955 1.465 ;
        RECT  0.100 1.205 0.310 1.705 ;
        END
        AntennaGateArea 0.3458 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.090 -0.130 11.480 0.130 ;
        RECT  10.830 -0.130 11.090 0.375 ;
        RECT  9.940 -0.130 10.830 0.130 ;
        RECT  9.680 -0.130 9.940 0.375 ;
        RECT  7.000 -0.130 9.680 0.130 ;
        RECT  6.400 -0.130 7.000 0.250 ;
        RECT  5.210 -0.130 6.400 0.130 ;
        RECT  4.610 -0.130 5.210 0.250 ;
        RECT  3.210 -0.130 4.610 0.130 ;
        RECT  2.270 -0.130 3.210 0.250 ;
        RECT  1.815 -0.130 2.270 0.130 ;
        RECT  1.215 -0.130 1.815 0.250 ;
        RECT  0.425 -0.130 1.215 0.130 ;
        RECT  0.165 -0.130 0.425 0.870 ;
        RECT  0.000 -0.130 0.165 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.505 2.740 11.480 3.000 ;
        RECT  10.245 2.305 10.505 3.000 ;
        RECT  8.765 2.740 10.245 3.000 ;
        RECT  8.265 2.195 8.765 3.000 ;
        RECT  5.210 2.740 8.265 3.000 ;
        RECT  4.610 2.620 5.210 3.000 ;
        RECT  3.210 2.740 4.610 3.000 ;
        RECT  2.270 2.620 3.210 3.000 ;
        RECT  1.325 2.740 2.270 3.000 ;
        RECT  1.065 1.985 1.325 3.000 ;
        RECT  0.000 2.740 1.065 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.780 1.045 10.880 1.205 ;
        RECT  10.620 1.045 10.780 1.675 ;
        RECT  9.845 1.515 10.620 1.675 ;
        RECT  10.065 1.005 10.345 1.305 ;
        RECT  9.045 1.005 10.065 1.165 ;
        RECT  9.245 1.345 9.845 1.675 ;
        RECT  8.590 1.515 9.245 1.675 ;
        RECT  8.930 1.005 9.045 1.335 ;
        RECT  8.770 0.310 8.930 1.335 ;
        RECT  7.375 0.310 8.770 0.470 ;
        RECT  8.430 0.650 8.590 1.945 ;
        RECT  7.710 0.650 8.430 0.810 ;
        RECT  8.240 1.685 8.430 1.945 ;
        RECT  8.050 1.035 8.250 1.195 ;
        RECT  7.890 1.035 8.050 2.560 ;
        RECT  5.980 2.400 7.890 2.560 ;
        RECT  7.550 0.650 7.710 2.220 ;
        RECT  6.750 2.060 7.550 2.220 ;
        RECT  7.215 0.310 7.375 0.590 ;
        RECT  7.185 0.785 7.370 1.865 ;
        RECT  5.980 0.430 7.215 0.590 ;
        RECT  6.930 0.785 7.185 0.945 ;
        RECT  6.930 1.705 7.185 1.865 ;
        RECT  6.750 1.215 6.890 1.475 ;
        RECT  6.590 0.810 6.750 2.220 ;
        RECT  4.000 0.810 6.590 0.970 ;
        RECT  5.810 1.705 6.590 1.865 ;
        RECT  3.795 1.235 6.410 1.495 ;
        RECT  5.380 0.310 5.980 0.590 ;
        RECT  5.380 2.280 5.980 2.560 ;
        RECT  5.550 1.705 5.810 1.995 ;
        RECT  4.210 1.705 5.550 1.865 ;
        RECT  4.430 0.430 5.380 0.590 ;
        RECT  4.430 2.280 5.380 2.440 ;
        RECT  4.235 0.310 4.430 0.590 ;
        RECT  4.170 2.280 4.430 2.560 ;
        RECT  4.170 0.310 4.235 0.565 ;
        RECT  4.050 1.705 4.210 1.965 ;
        RECT  3.490 0.405 4.170 0.565 ;
        RECT  1.885 2.280 4.170 2.440 ;
        RECT  3.635 0.765 3.795 2.005 ;
        RECT  3.540 0.765 3.635 1.025 ;
        RECT  3.540 1.685 3.635 2.005 ;
        RECT  3.330 0.405 3.490 0.590 ;
        RECT  3.360 1.210 3.455 1.470 ;
        RECT  3.200 0.815 3.360 2.030 ;
        RECT  1.420 0.430 3.330 0.590 ;
        RECT  2.550 0.815 3.200 0.975 ;
        RECT  2.115 1.870 3.200 2.030 ;
        RECT  1.725 0.770 1.885 2.440 ;
        RECT  1.615 0.770 1.725 0.995 ;
        RECT  1.605 1.825 1.725 2.440 ;
        RECT  1.420 1.245 1.535 1.505 ;
        RECT  1.260 0.430 1.420 1.805 ;
        RECT  0.935 0.710 1.260 0.870 ;
        RECT  0.785 1.645 1.260 1.805 ;
        RECT  0.675 0.610 0.935 0.870 ;
        RECT  0.525 1.645 0.785 2.325 ;
    END
END TLATNTSCAX6MTH

MACRO TLATNTSCAX8MTH
    CLASS CORE ;
    FOREIGN TLATNTSCAX8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 13.120 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SE
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.560 1.165 2.975 1.635 ;
        END
        AntennaGateArea 0.1222 ;
    END SE
    PIN ECK
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  12.610 0.435 12.990 2.125 ;
        RECT  9.920 0.435 12.610 0.775 ;
        RECT  12.230 1.740 12.610 2.125 ;
        RECT  12.155 1.740 12.230 2.465 ;
        RECT  11.850 1.865 12.155 2.465 ;
        RECT  10.550 1.865 11.850 2.125 ;
        RECT  10.170 1.865 10.550 2.465 ;
        END
        AntennaDiffArea 1.172 ;
    END ECK
    PIN E
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.065 1.120 2.380 1.680 ;
        END
        AntennaGateArea 0.1222 ;
    END E
    PIN CK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.205 0.955 1.465 ;
        RECT  0.100 1.205 0.310 1.705 ;
        END
        AntennaGateArea 0.4108 ;
    END CK
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.890 -0.130 13.120 0.130 ;
        RECT  11.950 -0.130 12.890 0.250 ;
        RECT  11.115 -0.130 11.950 0.130 ;
        RECT  10.515 -0.130 11.115 0.250 ;
        RECT  7.790 -0.130 10.515 0.130 ;
        RECT  7.190 -0.130 7.790 0.250 ;
        RECT  5.995 -0.130 7.190 0.130 ;
        RECT  5.395 -0.130 5.995 0.250 ;
        RECT  3.065 -0.130 5.395 0.130 ;
        RECT  2.125 -0.130 3.065 0.250 ;
        RECT  1.475 -0.130 2.125 0.130 ;
        RECT  1.215 -0.130 1.475 0.250 ;
        RECT  0.425 -0.130 1.215 0.130 ;
        RECT  0.165 -0.130 0.425 0.975 ;
        RECT  0.000 -0.130 0.165 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  12.995 2.740 13.120 3.000 ;
        RECT  12.735 2.305 12.995 3.000 ;
        RECT  11.320 2.740 12.735 3.000 ;
        RECT  11.060 2.305 11.320 3.000 ;
        RECT  9.570 2.740 11.060 3.000 ;
        RECT  9.070 2.195 9.570 3.000 ;
        RECT  5.995 2.740 9.070 3.000 ;
        RECT  5.395 2.620 5.995 3.000 ;
        RECT  4.075 2.740 5.395 3.000 ;
        RECT  3.135 2.620 4.075 3.000 ;
        RECT  2.605 2.740 3.135 3.000 ;
        RECT  1.665 2.620 2.605 3.000 ;
        RECT  1.325 2.740 1.665 3.000 ;
        RECT  1.065 1.985 1.325 3.000 ;
        RECT  0.000 2.740 1.065 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  12.270 0.965 12.430 1.225 ;
        RECT  11.480 0.995 12.270 1.155 ;
        RECT  11.975 1.335 12.000 1.585 ;
        RECT  11.740 1.335 11.975 1.685 ;
        RECT  10.660 1.525 11.740 1.685 ;
        RECT  10.880 0.995 11.480 1.345 ;
        RECT  9.785 0.995 10.880 1.155 ;
        RECT  10.060 1.335 10.660 1.685 ;
        RECT  9.345 1.525 10.060 1.685 ;
        RECT  9.685 0.995 9.785 1.345 ;
        RECT  9.525 0.310 9.685 1.345 ;
        RECT  8.180 0.310 9.525 0.470 ;
        RECT  9.185 0.650 9.345 1.945 ;
        RECT  8.515 0.650 9.185 0.810 ;
        RECT  9.045 1.685 9.185 1.945 ;
        RECT  8.855 1.005 9.005 1.265 ;
        RECT  8.695 1.005 8.855 2.560 ;
        RECT  6.770 2.400 8.695 2.560 ;
        RECT  8.355 0.650 8.515 2.220 ;
        RECT  7.555 2.060 8.355 2.220 ;
        RECT  8.020 0.310 8.180 0.590 ;
        RECT  7.990 0.785 8.175 1.865 ;
        RECT  6.770 0.430 8.020 0.590 ;
        RECT  7.735 0.785 7.990 0.945 ;
        RECT  7.735 1.705 7.990 1.865 ;
        RECT  7.555 1.215 7.695 1.475 ;
        RECT  7.395 0.770 7.555 2.220 ;
        RECT  4.790 0.770 7.395 0.930 ;
        RECT  4.790 1.755 7.395 1.915 ;
        RECT  4.300 1.235 7.200 1.495 ;
        RECT  6.170 0.310 6.770 0.590 ;
        RECT  6.170 2.100 6.770 2.560 ;
        RECT  5.220 0.430 6.170 0.590 ;
        RECT  5.220 2.100 6.170 2.260 ;
        RECT  4.780 0.310 5.220 0.590 ;
        RECT  4.620 2.100 5.220 2.560 ;
        RECT  4.620 0.310 4.780 0.565 ;
        RECT  3.365 0.405 4.620 0.565 ;
        RECT  1.885 2.210 4.620 2.370 ;
        RECT  4.140 0.865 4.300 1.845 ;
        RECT  3.700 0.865 4.140 1.025 ;
        RECT  3.700 1.685 4.140 1.845 ;
        RECT  3.360 1.210 3.920 1.470 ;
        RECT  3.540 0.765 3.700 1.025 ;
        RECT  3.540 1.685 3.700 1.945 ;
        RECT  3.205 0.405 3.365 0.590 ;
        RECT  3.200 0.775 3.360 2.030 ;
        RECT  1.420 0.430 3.205 0.590 ;
        RECT  2.550 0.775 3.200 0.935 ;
        RECT  2.115 1.870 3.200 2.030 ;
        RECT  1.725 0.815 1.885 2.370 ;
        RECT  1.615 0.815 1.725 0.975 ;
        RECT  1.605 1.865 1.725 2.370 ;
        RECT  1.420 1.245 1.535 1.505 ;
        RECT  1.260 0.430 1.420 1.805 ;
        RECT  0.935 0.815 1.260 0.975 ;
        RECT  0.785 1.645 1.260 1.805 ;
        RECT  0.675 0.375 0.935 0.975 ;
        RECT  0.525 1.645 0.785 2.405 ;
    END
END TLATNTSCAX8MTH

MACRO TLATNX1MTH
    CLASS CORE ;
    FOREIGN TLATNX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 0.735 5.640 2.020 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.595 1.290 4.820 1.580 ;
        RECT  4.335 0.815 4.595 2.015 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.395 1.790 ;
        END
        AntennaGateArea 0.0741 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.615 0.880 2.005 1.365 ;
        END
        AntennaGateArea 0.1534 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.135 -0.130 5.740 0.130 ;
        RECT  4.875 -0.130 5.135 0.295 ;
        RECT  3.515 -0.130 4.875 0.130 ;
        RECT  3.255 -0.130 3.515 0.310 ;
        RECT  1.805 -0.130 3.255 0.130 ;
        RECT  1.545 -0.130 1.805 0.360 ;
        RECT  0.385 -0.130 1.545 0.130 ;
        RECT  0.125 -0.130 0.385 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.105 2.740 5.740 3.000 ;
        RECT  4.845 1.760 5.105 3.000 ;
        RECT  3.595 2.740 4.845 3.000 ;
        RECT  3.335 2.345 3.595 3.000 ;
        RECT  1.805 2.740 3.335 3.000 ;
        RECT  1.545 2.615 1.805 3.000 ;
        RECT  0.385 2.740 1.545 3.000 ;
        RECT  0.125 2.285 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.040 0.475 5.200 1.495 ;
        RECT  4.035 0.475 5.040 0.635 ;
        RECT  3.875 0.475 4.035 2.125 ;
        RECT  3.405 1.440 3.875 1.600 ;
        RECT  3.535 0.960 3.695 1.220 ;
        RECT  2.870 1.060 3.535 1.220 ;
        RECT  3.145 1.440 3.405 1.700 ;
        RECT  2.240 0.310 2.915 0.470 ;
        RECT  2.725 2.400 2.915 2.560 ;
        RECT  2.710 0.715 2.870 2.075 ;
        RECT  2.565 2.275 2.725 2.560 ;
        RECT  2.435 0.715 2.710 0.975 ;
        RECT  2.435 1.915 2.710 2.075 ;
        RECT  0.765 2.275 2.565 2.435 ;
        RECT  1.275 1.545 2.485 1.705 ;
        RECT  2.080 0.310 2.240 0.700 ;
        RECT  1.275 0.540 2.080 0.700 ;
        RECT  1.115 0.540 1.275 2.055 ;
        RECT  0.765 1.220 0.905 1.480 ;
        RECT  0.605 0.765 0.765 2.435 ;
    END
END TLATNX1MTH

MACRO TLATNX2MTH
    CLASS CORE ;
    FOREIGN TLATNX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 0.385 5.640 2.415 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 0.815 4.595 2.415 ;
        RECT  4.275 0.815 4.335 0.975 ;
        RECT  4.200 1.285 4.335 1.580 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.395 1.790 ;
        END
        AntennaGateArea 0.0897 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 0.855 1.995 1.345 ;
        END
        AntennaGateArea 0.1833 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 -0.130 5.740 0.130 ;
        RECT  4.815 -0.130 5.075 0.290 ;
        RECT  3.455 -0.130 4.815 0.130 ;
        RECT  3.195 -0.130 3.455 0.340 ;
        RECT  1.795 -0.130 3.195 0.130 ;
        RECT  1.195 -0.130 1.795 0.300 ;
        RECT  0.725 -0.130 1.195 0.130 ;
        RECT  0.125 -0.130 0.725 0.300 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.105 2.740 5.740 3.000 ;
        RECT  4.845 1.815 5.105 3.000 ;
        RECT  3.530 2.740 4.845 3.000 ;
        RECT  3.270 2.240 3.530 3.000 ;
        RECT  1.835 2.740 3.270 3.000 ;
        RECT  0.895 2.620 1.835 3.000 ;
        RECT  0.385 2.740 0.895 3.000 ;
        RECT  0.125 2.315 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.040 0.475 5.200 1.480 ;
        RECT  4.020 0.475 5.040 0.635 ;
        RECT  3.860 0.475 4.020 2.110 ;
        RECT  3.805 0.475 3.860 0.810 ;
        RECT  3.370 1.420 3.860 1.580 ;
        RECT  3.520 0.940 3.680 1.200 ;
        RECT  3.030 1.040 3.520 1.200 ;
        RECT  3.210 1.420 3.370 1.680 ;
        RECT  2.180 2.400 3.075 2.560 ;
        RECT  2.870 0.815 3.030 2.120 ;
        RECT  2.185 0.310 2.905 0.470 ;
        RECT  2.645 0.815 2.870 0.975 ;
        RECT  2.445 1.960 2.870 2.120 ;
        RECT  2.385 0.715 2.645 0.975 ;
        RECT  2.275 1.500 2.535 1.690 ;
        RECT  1.245 1.530 2.275 1.690 ;
        RECT  2.025 0.310 2.185 0.670 ;
        RECT  2.020 2.280 2.180 2.560 ;
        RECT  1.245 0.510 2.025 0.670 ;
        RECT  0.735 2.280 2.020 2.440 ;
        RECT  1.085 0.510 1.245 2.100 ;
        RECT  0.735 1.220 0.875 1.480 ;
        RECT  0.575 0.760 0.735 2.440 ;
    END
END TLATNX2MTH

MACRO TLATNX4MTH
    CLASS CORE ;
    FOREIGN TLATNX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.945 1.290 6.050 1.580 ;
        RECT  5.765 0.385 5.945 2.410 ;
        RECT  5.665 0.385 5.765 0.985 ;
        RECT  5.665 1.810 5.765 2.410 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 0.810 4.985 2.410 ;
        RECT  4.605 1.290 4.725 1.580 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN GN
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.505 1.595 ;
        END
        AntennaGateArea 0.1677 ;
    END GN
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 0.855 2.095 1.350 ;
        END
        AntennaGateArea 0.182 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.985 ;
        RECT  4.445 -0.130 6.175 0.130 ;
        RECT  4.185 -0.130 4.445 0.280 ;
        RECT  3.515 -0.130 4.185 0.130 ;
        RECT  3.255 -0.130 3.515 0.300 ;
        RECT  1.855 -0.130 3.255 0.130 ;
        RECT  1.595 -0.130 1.855 0.250 ;
        RECT  0.385 -0.130 1.595 0.130 ;
        RECT  0.125 -0.130 0.385 0.880 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.805 6.435 3.000 ;
        RECT  4.445 2.740 6.175 3.000 ;
        RECT  4.185 2.325 4.445 3.000 ;
        RECT  3.465 2.740 4.185 3.000 ;
        RECT  3.205 2.275 3.465 3.000 ;
        RECT  1.825 2.740 3.205 3.000 ;
        RECT  1.565 2.530 1.825 3.000 ;
        RECT  0.385 2.740 1.565 3.000 ;
        RECT  0.125 1.775 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.485 1.200 5.585 1.460 ;
        RECT  5.325 0.460 5.485 1.460 ;
        RECT  4.175 0.460 5.325 0.620 ;
        RECT  4.015 0.460 4.175 2.125 ;
        RECT  3.795 0.685 4.015 0.945 ;
        RECT  3.745 1.545 4.015 2.125 ;
        RECT  2.875 1.185 3.835 1.345 ;
        RECT  3.095 1.545 3.745 1.705 ;
        RECT  2.220 0.310 2.965 0.470 ;
        RECT  2.215 2.400 2.960 2.560 ;
        RECT  2.715 0.655 2.875 2.030 ;
        RECT  2.470 0.655 2.715 0.915 ;
        RECT  2.675 1.870 2.715 2.030 ;
        RECT  2.415 1.870 2.675 2.130 ;
        RECT  1.355 1.530 2.535 1.690 ;
        RECT  2.060 0.310 2.220 0.590 ;
        RECT  2.055 2.190 2.215 2.560 ;
        RECT  1.355 0.430 2.060 0.590 ;
        RECT  0.845 2.190 2.055 2.350 ;
        RECT  1.195 0.430 1.355 2.010 ;
        RECT  0.845 1.240 0.985 1.500 ;
        RECT  0.685 0.620 0.845 2.350 ;
    END
END TLATNX4MTH

MACRO TLATSRX1MTH
    CLASS CORE ;
    FOREIGN TLATSRX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.140 0.515 1.605 ;
        END
        AntennaGateArea 0.0897 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.595 0.920 2.810 1.470 ;
        RECT  2.520 0.920 2.595 1.130 ;
        END
        AntennaGateArea 0.1456 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.350 0.705 8.510 2.000 ;
        RECT  8.275 0.705 8.350 0.965 ;
        RECT  8.270 1.700 8.350 2.000 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.530 1.265 7.690 1.580 ;
        RECT  7.530 0.815 7.555 0.975 ;
        RECT  7.370 0.815 7.530 1.895 ;
        RECT  7.295 0.815 7.370 0.975 ;
        RECT  7.270 1.735 7.370 1.895 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.820 1.190 5.155 1.505 ;
        RECT  4.610 0.880 4.820 1.505 ;
        END
        AntennaGateArea 0.0793 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.885 1.295 2.400 1.540 ;
        END
        AntennaGateArea 0.1183 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  8.435 -0.130 8.610 0.130 ;
        RECT  7.835 -0.130 8.435 0.285 ;
        RECT  7.535 -0.130 7.835 0.130 ;
        RECT  6.935 -0.130 7.535 0.285 ;
        RECT  6.590 -0.130 6.935 0.130 ;
        RECT  5.990 -0.130 6.590 0.275 ;
        RECT  5.770 -0.130 5.990 0.130 ;
        RECT  4.830 -0.130 5.770 0.275 ;
        RECT  2.305 -0.130 4.830 0.130 ;
        RECT  1.805 -0.130 2.305 0.365 ;
        RECT  0.385 -0.130 1.805 0.130 ;
        RECT  0.125 -0.130 0.385 0.475 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.940 2.740 8.610 3.000 ;
        RECT  7.340 2.620 7.940 3.000 ;
        RECT  0.440 2.740 7.340 3.000 ;
        RECT  0.180 2.315 0.440 3.000 ;
        RECT  0.000 2.740 0.180 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.090 1.150 8.155 1.410 ;
        RECT  7.930 0.470 8.090 2.415 ;
        RECT  6.995 0.470 7.930 0.630 ;
        RECT  6.970 2.255 7.930 2.415 ;
        RECT  6.630 1.200 7.190 1.460 ;
        RECT  6.835 0.470 6.995 1.005 ;
        RECT  6.810 1.700 6.970 2.560 ;
        RECT  4.255 2.400 6.810 2.560 ;
        RECT  6.590 1.200 6.630 2.220 ;
        RECT  6.470 1.255 6.590 2.220 ;
        RECT  1.365 2.060 6.470 2.220 ;
        RECT  6.130 0.850 6.290 1.880 ;
        RECT  6.005 0.850 6.130 1.010 ;
        RECT  5.695 1.720 6.130 1.880 ;
        RECT  5.845 0.455 6.005 1.010 ;
        RECT  5.495 1.220 5.950 1.480 ;
        RECT  5.045 0.455 5.845 0.615 ;
        RECT  5.495 0.795 5.545 0.955 ;
        RECT  5.335 0.795 5.495 1.880 ;
        RECT  5.285 0.795 5.335 0.955 ;
        RECT  3.150 1.720 5.335 1.880 ;
        RECT  4.885 0.455 5.045 0.700 ;
        RECT  4.420 0.540 4.885 0.700 ;
        RECT  4.260 0.540 4.420 1.540 ;
        RECT  3.600 1.380 4.260 1.540 ;
        RECT  3.820 1.010 4.080 1.200 ;
        RECT  0.855 2.400 4.035 2.560 ;
        RECT  3.275 0.580 3.875 0.830 ;
        RECT  3.150 1.010 3.820 1.170 ;
        RECT  3.340 1.350 3.600 1.540 ;
        RECT  2.340 0.580 3.275 0.740 ;
        RECT  2.990 1.010 3.150 1.880 ;
        RECT  1.705 1.720 2.990 1.880 ;
        RECT  2.180 0.580 2.340 0.915 ;
        RECT  1.195 0.755 2.180 0.915 ;
        RECT  1.545 1.315 1.705 1.880 ;
        RECT  0.855 0.375 1.625 0.535 ;
        RECT  1.375 1.315 1.545 1.625 ;
        RECT  1.205 1.815 1.365 2.220 ;
        RECT  1.195 1.815 1.205 1.975 ;
        RECT  1.035 0.755 1.195 1.975 ;
        RECT  0.695 0.375 0.855 2.560 ;
    END
END TLATSRX1MTH

MACRO TLATSRX2MTH
    CLASS CORE ;
    FOREIGN TLATSRX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.610 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 0.880 0.395 1.495 ;
        END
        AntennaGateArea 0.13 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.310 2.855 1.470 ;
        RECT  2.560 0.880 2.780 1.470 ;
        END
        AntennaGateArea 0.182 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.350 0.355 8.510 2.465 ;
        RECT  8.275 0.355 8.350 0.955 ;
        RECT  8.270 1.700 8.350 2.465 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 1.285 7.750 1.580 ;
        RECT  7.375 0.815 7.535 1.895 ;
        RECT  7.275 0.815 7.375 0.975 ;
        RECT  7.145 1.735 7.375 1.895 ;
        END
        AntennaDiffArea 0.467 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.780 1.245 5.270 1.540 ;
        END
        AntennaGateArea 0.0858 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 0.880 2.375 1.455 ;
        END
        AntennaGateArea 0.1651 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.070 -0.130 8.610 0.130 ;
        RECT  6.130 -0.130 7.070 0.290 ;
        RECT  2.315 -0.130 6.130 0.130 ;
        RECT  1.715 -0.130 2.315 0.300 ;
        RECT  0.385 -0.130 1.715 0.130 ;
        RECT  0.125 -0.130 0.385 0.325 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 2.740 8.610 3.000 ;
        RECT  7.685 2.415 7.945 3.000 ;
        RECT  0.385 2.740 7.685 3.000 ;
        RECT  0.125 2.485 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.090 1.140 8.155 1.400 ;
        RECT  7.930 0.470 8.090 2.235 ;
        RECT  7.025 0.470 7.930 0.630 ;
        RECT  6.955 2.075 7.930 2.235 ;
        RECT  6.590 1.220 7.195 1.480 ;
        RECT  6.865 0.470 7.025 0.840 ;
        RECT  6.795 2.075 6.955 2.560 ;
        RECT  6.765 0.680 6.865 0.840 ;
        RECT  4.255 2.400 6.795 2.560 ;
        RECT  6.430 1.220 6.590 2.220 ;
        RECT  1.855 2.060 6.430 2.220 ;
        RECT  6.090 0.730 6.250 1.780 ;
        RECT  6.005 0.730 6.090 0.890 ;
        RECT  5.950 1.620 6.090 1.780 ;
        RECT  5.950 0.630 6.005 0.890 ;
        RECT  5.790 0.410 5.950 0.890 ;
        RECT  5.790 1.620 5.950 1.880 ;
        RECT  5.610 1.180 5.910 1.440 ;
        RECT  5.100 0.410 5.790 0.570 ;
        RECT  5.450 0.750 5.610 1.880 ;
        RECT  5.285 0.750 5.450 0.910 ;
        RECT  3.200 1.720 5.450 1.880 ;
        RECT  4.910 0.410 5.100 0.620 ;
        RECT  4.475 0.460 4.910 0.620 ;
        RECT  4.315 0.460 4.475 1.540 ;
        RECT  3.655 1.380 4.315 1.540 ;
        RECT  3.875 1.010 4.135 1.200 ;
        RECT  0.735 2.400 4.050 2.560 ;
        RECT  3.275 0.540 3.875 0.830 ;
        RECT  3.200 1.010 3.875 1.170 ;
        RECT  3.395 1.350 3.655 1.540 ;
        RECT  1.660 0.540 3.275 0.700 ;
        RECT  3.040 1.010 3.200 1.880 ;
        RECT  2.290 1.720 3.040 1.880 ;
        RECT  2.130 1.645 2.290 1.880 ;
        RECT  1.415 1.645 2.130 1.805 ;
        RECT  1.695 2.005 1.855 2.220 ;
        RECT  1.075 2.005 1.695 2.165 ;
        RECT  1.500 0.540 1.660 0.865 ;
        RECT  1.075 0.705 1.500 0.865 ;
        RECT  1.255 1.315 1.415 1.805 ;
        RECT  0.735 0.335 1.155 0.495 ;
        RECT  0.915 0.705 1.075 2.165 ;
        RECT  0.575 0.335 0.735 2.560 ;
    END
END TLATSRX2MTH

MACRO TLATSRX4MTH
    CLASS CORE ;
    FOREIGN TLATSRX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.840 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN SN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.235 0.395 1.660 ;
        END
        AntennaGateArea 0.1638 ;
    END SN
    PIN RN
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.780 1.310 2.855 1.470 ;
        RECT  2.560 0.880 2.780 1.470 ;
        END
        AntennaGateArea 0.182 ;
    END RN
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.235 1.290 9.330 1.580 ;
        RECT  9.055 0.355 9.235 2.390 ;
        RECT  8.945 0.355 9.055 0.955 ;
        RECT  8.945 1.790 9.055 2.390 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.965 0.360 8.185 0.960 ;
        RECT  7.805 0.360 7.965 2.065 ;
        RECT  7.480 1.675 7.805 2.065 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  4.735 1.190 5.270 1.540 ;
        END
        AntennaGateArea 0.1391 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.115 0.880 2.375 1.455 ;
        END
        AntennaGateArea 0.1651 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.715 -0.130 9.840 0.130 ;
        RECT  9.455 -0.130 9.715 0.955 ;
        RECT  8.695 -0.130 9.455 0.130 ;
        RECT  8.435 -0.130 8.695 0.955 ;
        RECT  7.625 -0.130 8.435 0.130 ;
        RECT  7.465 -0.130 7.625 1.025 ;
        RECT  6.625 -0.130 7.465 0.130 ;
        RECT  6.365 -0.130 6.625 0.670 ;
        RECT  5.025 -0.130 6.365 0.130 ;
        RECT  4.765 -0.130 5.025 0.280 ;
        RECT  2.420 -0.130 4.765 0.130 ;
        RECT  1.820 -0.130 2.420 0.355 ;
        RECT  0.385 -0.130 1.820 0.130 ;
        RECT  0.125 -0.130 0.385 0.855 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.715 2.740 9.840 3.000 ;
        RECT  9.455 1.790 9.715 3.000 ;
        RECT  8.645 2.740 9.455 3.000 ;
        RECT  8.485 1.790 8.645 3.000 ;
        RECT  8.305 2.595 8.485 3.000 ;
        RECT  7.475 2.740 8.305 3.000 ;
        RECT  7.215 2.595 7.475 3.000 ;
        RECT  0.385 2.740 7.215 3.000 ;
        RECT  0.125 2.620 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.305 1.140 8.875 1.400 ;
        RECT  8.145 1.140 8.305 2.415 ;
        RECT  7.045 2.255 8.145 2.415 ;
        RECT  7.045 0.650 7.115 0.910 ;
        RECT  7.025 0.650 7.045 2.415 ;
        RECT  6.885 0.650 7.025 2.560 ;
        RECT  6.840 1.845 6.885 2.560 ;
        RECT  4.255 2.400 6.840 2.560 ;
        RECT  6.630 1.185 6.705 1.445 ;
        RECT  6.470 1.185 6.630 2.220 ;
        RECT  1.855 2.060 6.470 2.220 ;
        RECT  6.130 0.850 6.290 1.880 ;
        RECT  6.035 0.850 6.130 1.010 ;
        RECT  5.790 1.720 6.130 1.880 ;
        RECT  5.875 0.460 6.035 1.010 ;
        RECT  5.610 1.220 5.950 1.480 ;
        RECT  5.125 0.460 5.875 0.620 ;
        RECT  5.450 0.800 5.610 1.880 ;
        RECT  5.315 0.800 5.450 0.960 ;
        RECT  3.200 1.720 5.450 1.880 ;
        RECT  4.965 0.460 5.125 0.885 ;
        RECT  4.475 0.725 4.965 0.885 ;
        RECT  4.315 0.725 4.475 1.540 ;
        RECT  3.655 1.380 4.315 1.540 ;
        RECT  3.875 1.010 4.135 1.200 ;
        RECT  0.735 2.400 4.050 2.560 ;
        RECT  3.275 0.540 3.875 0.830 ;
        RECT  3.200 1.010 3.875 1.170 ;
        RECT  3.395 1.350 3.655 1.540 ;
        RECT  1.660 0.540 3.275 0.700 ;
        RECT  3.040 1.010 3.200 1.880 ;
        RECT  2.290 1.720 3.040 1.880 ;
        RECT  2.130 1.645 2.290 1.880 ;
        RECT  1.535 1.645 2.130 1.805 ;
        RECT  1.695 2.005 1.855 2.220 ;
        RECT  1.195 2.005 1.695 2.165 ;
        RECT  1.500 0.540 1.660 0.865 ;
        RECT  1.375 1.315 1.535 1.805 ;
        RECT  1.195 0.705 1.500 0.865 ;
        RECT  0.845 0.335 1.265 0.495 ;
        RECT  1.035 0.705 1.195 2.165 ;
        RECT  0.735 0.335 0.845 0.975 ;
        RECT  0.575 0.335 0.735 2.560 ;
    END
END TLATSRX4MTH

MACRO TLATX1MTH
    CLASS CORE ;
    FOREIGN TLATX1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 0.735 5.640 2.145 ;
        END
        AntennaDiffArea 0.333 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 0.815 4.595 2.080 ;
        RECT  4.200 0.815 4.335 1.580 ;
        END
        AntennaDiffArea 0.333 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.395 1.790 ;
        END
        AntennaGateArea 0.0663 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.735 0.855 1.975 1.650 ;
        END
        AntennaGateArea 0.1534 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 -0.130 5.740 0.130 ;
        RECT  4.815 -0.130 5.075 0.250 ;
        RECT  3.455 -0.130 4.815 0.130 ;
        RECT  3.195 -0.130 3.455 0.340 ;
        RECT  1.795 -0.130 3.195 0.130 ;
        RECT  1.535 -0.130 1.795 0.250 ;
        RECT  0.385 -0.130 1.535 0.130 ;
        RECT  0.125 -0.130 0.385 0.465 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.105 2.740 5.740 3.000 ;
        RECT  4.845 1.970 5.105 3.000 ;
        RECT  3.570 2.740 4.845 3.000 ;
        RECT  3.310 2.525 3.570 3.000 ;
        RECT  1.820 2.740 3.310 3.000 ;
        RECT  1.560 2.235 1.820 3.000 ;
        RECT  0.385 2.740 1.560 3.000 ;
        RECT  0.125 2.315 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.040 0.475 5.200 1.485 ;
        RECT  4.020 0.475 5.040 0.635 ;
        RECT  4.020 2.045 4.085 2.305 ;
        RECT  3.860 0.475 4.020 2.305 ;
        RECT  3.815 0.475 3.860 0.735 ;
        RECT  3.335 1.395 3.860 1.555 ;
        RECT  3.520 0.915 3.680 1.175 ;
        RECT  2.995 1.015 3.520 1.175 ;
        RECT  3.175 1.395 3.335 1.655 ;
        RECT  2.835 0.785 2.995 2.005 ;
        RECT  2.315 2.395 2.935 2.555 ;
        RECT  2.180 0.310 2.905 0.470 ;
        RECT  2.645 0.785 2.835 0.945 ;
        RECT  2.655 1.845 2.835 2.005 ;
        RECT  2.495 1.845 2.655 2.105 ;
        RECT  2.385 0.685 2.645 0.945 ;
        RECT  2.315 1.125 2.510 1.285 ;
        RECT  2.155 1.125 2.315 2.555 ;
        RECT  2.020 0.310 2.180 0.590 ;
        RECT  1.275 1.855 2.155 2.015 ;
        RECT  0.765 0.430 2.020 0.590 ;
        RECT  1.275 0.770 1.325 0.930 ;
        RECT  1.115 0.770 1.275 2.015 ;
        RECT  1.065 0.770 1.115 0.930 ;
        RECT  0.765 1.220 0.875 1.480 ;
        RECT  0.605 0.430 0.765 1.980 ;
    END
END TLATX1MTH

MACRO TLATX2MTH
    CLASS CORE ;
    FOREIGN TLATX2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.380 0.375 5.640 2.405 ;
        END
        AntennaDiffArea 0.537 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.335 0.815 4.595 2.405 ;
        RECT  4.200 0.815 4.335 1.580 ;
        END
        AntennaDiffArea 0.537 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.395 1.790 ;
        END
        AntennaGateArea 0.0871 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.565 0.855 1.950 1.395 ;
        END
        AntennaGateArea 0.1885 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.075 -0.130 5.740 0.130 ;
        RECT  4.815 -0.130 5.075 0.250 ;
        RECT  3.455 -0.130 4.815 0.130 ;
        RECT  3.195 -0.130 3.455 0.340 ;
        RECT  1.795 -0.130 3.195 0.130 ;
        RECT  1.535 -0.130 1.795 0.250 ;
        RECT  0.385 -0.130 1.535 0.130 ;
        RECT  0.125 -0.130 0.385 0.465 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.105 2.740 5.740 3.000 ;
        RECT  4.845 1.805 5.105 3.000 ;
        RECT  3.545 2.740 4.845 3.000 ;
        RECT  3.285 2.455 3.545 3.000 ;
        RECT  1.795 2.740 3.285 3.000 ;
        RECT  1.535 2.235 1.795 3.000 ;
        RECT  0.385 2.740 1.535 3.000 ;
        RECT  0.125 2.315 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.040 0.475 5.200 1.485 ;
        RECT  4.020 0.475 5.040 0.635 ;
        RECT  4.020 1.850 4.085 2.110 ;
        RECT  3.860 0.475 4.020 2.110 ;
        RECT  3.815 0.475 3.860 0.735 ;
        RECT  3.380 1.420 3.860 1.580 ;
        RECT  3.520 0.940 3.680 1.200 ;
        RECT  3.030 1.040 3.520 1.200 ;
        RECT  3.220 1.420 3.380 1.680 ;
        RECT  2.870 0.785 3.030 2.005 ;
        RECT  2.180 0.310 2.905 0.470 ;
        RECT  2.315 2.325 2.905 2.485 ;
        RECT  2.645 0.785 2.870 0.945 ;
        RECT  2.655 1.845 2.870 2.005 ;
        RECT  2.495 1.845 2.655 2.105 ;
        RECT  2.385 0.685 2.645 0.945 ;
        RECT  2.315 1.125 2.475 1.285 ;
        RECT  2.155 1.125 2.315 2.485 ;
        RECT  2.020 0.310 2.180 0.590 ;
        RECT  1.245 1.855 2.155 2.015 ;
        RECT  0.735 0.430 2.020 0.590 ;
        RECT  1.245 0.815 1.295 0.975 ;
        RECT  1.085 0.815 1.245 2.015 ;
        RECT  1.035 0.815 1.085 0.975 ;
        RECT  0.735 1.220 0.875 1.480 ;
        RECT  0.575 0.430 0.735 1.980 ;
    END
END TLATX2MTH

MACRO TLATX4MTH
    CLASS CORE ;
    FOREIGN TLATX4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.560 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN QN
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.925 1.290 6.050 1.580 ;
        RECT  5.765 0.390 5.925 2.415 ;
        RECT  5.665 0.390 5.765 0.990 ;
        RECT  5.665 1.815 5.765 2.415 ;
        END
        AntennaDiffArea 0.6 ;
    END QN
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.725 0.800 4.985 2.415 ;
        RECT  4.605 1.290 4.725 1.580 ;
        END
        AntennaDiffArea 0.6 ;
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.505 1.595 ;
        END
        AntennaGateArea 0.1677 ;
    END G
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.665 0.855 2.005 1.405 ;
        END
        AntennaGateArea 0.182 ;
    END D
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 -0.130 6.560 0.130 ;
        RECT  6.175 -0.130 6.435 0.985 ;
        RECT  4.445 -0.130 6.175 0.130 ;
        RECT  4.185 -0.130 4.445 0.280 ;
        RECT  3.515 -0.130 4.185 0.130 ;
        RECT  3.255 -0.130 3.515 0.360 ;
        RECT  1.855 -0.130 3.255 0.130 ;
        RECT  1.595 -0.130 1.855 0.295 ;
        RECT  0.385 -0.130 1.595 0.130 ;
        RECT  0.125 -0.130 0.385 0.880 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  6.435 2.740 6.560 3.000 ;
        RECT  6.175 1.815 6.435 3.000 ;
        RECT  4.445 2.740 6.175 3.000 ;
        RECT  4.185 2.565 4.445 3.000 ;
        RECT  3.465 2.740 4.185 3.000 ;
        RECT  3.205 2.535 3.465 3.000 ;
        RECT  1.805 2.740 3.205 3.000 ;
        RECT  1.545 2.485 1.805 3.000 ;
        RECT  0.385 2.740 1.545 3.000 ;
        RECT  0.125 1.790 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.485 1.200 5.585 1.460 ;
        RECT  5.325 0.460 5.485 1.460 ;
        RECT  4.175 0.460 5.325 0.620 ;
        RECT  4.015 0.460 4.175 2.125 ;
        RECT  3.795 0.685 4.015 0.945 ;
        RECT  3.745 1.545 4.015 2.125 ;
        RECT  2.875 1.185 3.835 1.345 ;
        RECT  3.095 1.545 3.745 1.705 ;
        RECT  2.220 0.310 2.965 0.470 ;
        RECT  2.215 2.400 2.915 2.560 ;
        RECT  2.715 0.650 2.875 2.220 ;
        RECT  2.445 0.650 2.715 0.915 ;
        RECT  2.445 1.960 2.715 2.220 ;
        RECT  2.435 1.185 2.535 1.345 ;
        RECT  2.275 1.185 2.435 1.745 ;
        RECT  2.215 1.585 2.275 1.745 ;
        RECT  2.060 0.310 2.220 0.635 ;
        RECT  2.055 1.585 2.215 2.560 ;
        RECT  0.845 0.475 2.060 0.635 ;
        RECT  1.355 1.930 2.055 2.090 ;
        RECT  1.355 0.815 1.405 0.975 ;
        RECT  1.195 0.815 1.355 2.090 ;
        RECT  1.145 0.815 1.195 0.975 ;
        RECT  0.845 1.220 1.015 1.480 ;
        RECT  0.685 0.475 0.845 2.355 ;
    END
END TLATX4MTH

MACRO XNOR2X1MTH
    CLASS CORE ;
    FOREIGN XNOR2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 1.290 3.590 1.580 ;
        RECT  3.365 1.290 3.465 1.945 ;
        RECT  3.205 0.765 3.365 1.945 ;
        RECT  3.095 0.765 3.205 1.025 ;
        END
        AntennaDiffArea 0.258 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.195 0.505 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.645 1.215 2.065 1.580 ;
        END
        AntennaGateArea 0.1417 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.260 -0.130 4.100 0.130 ;
        RECT  2.320 -0.130 3.260 0.250 ;
        RECT  1.605 -0.130 2.320 0.130 ;
        RECT  0.665 -0.130 1.605 0.250 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.875 2.740 4.100 3.000 ;
        RECT  0.935 2.570 1.875 3.000 ;
        RECT  0.605 2.740 0.935 3.000 ;
        RECT  0.345 2.555 0.605 3.000 ;
        RECT  0.000 2.740 0.345 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.770 0.765 3.930 2.285 ;
        RECT  3.605 0.765 3.770 1.025 ;
        RECT  3.715 1.730 3.770 2.285 ;
        RECT  0.930 2.125 3.715 2.285 ;
        RECT  2.915 1.685 2.955 1.945 ;
        RECT  2.755 0.475 2.915 1.945 ;
        RECT  2.585 0.475 2.755 1.025 ;
        RECT  2.695 1.685 2.755 1.945 ;
        RECT  1.325 0.475 2.585 0.635 ;
        RECT  2.405 1.255 2.575 1.515 ;
        RECT  2.405 1.760 2.445 1.920 ;
        RECT  2.245 0.815 2.405 1.920 ;
        RECT  2.075 0.815 2.245 0.975 ;
        RECT  2.185 1.760 2.245 1.920 ;
        RECT  1.325 1.685 1.375 1.945 ;
        RECT  1.165 0.475 1.325 1.945 ;
        RECT  1.115 1.685 1.165 1.945 ;
        RECT  0.930 1.225 0.985 1.485 ;
        RECT  0.770 0.830 0.930 2.285 ;
        RECT  0.385 0.830 0.770 0.990 ;
        RECT  0.385 1.760 0.770 1.920 ;
        RECT  0.125 0.730 0.385 0.990 ;
        RECT  0.125 1.760 0.385 2.020 ;
    END
END XNOR2X1MTH

MACRO XNOR2X2MTH
    CLASS CORE ;
    FOREIGN XNOR2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.345 1.290 3.590 1.580 ;
        RECT  3.345 1.845 3.465 2.005 ;
        RECT  3.345 0.565 3.395 0.825 ;
        RECT  3.185 0.565 3.345 2.005 ;
        RECT  3.135 0.565 3.185 0.825 ;
        END
        AntennaDiffArea 0.516 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.555 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.635 1.215 2.090 1.580 ;
        END
        AntennaGateArea 0.2522 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 -0.130 4.100 0.130 ;
        RECT  1.715 -0.130 1.975 0.285 ;
        RECT  0.925 -0.130 1.715 0.130 ;
        RECT  0.665 -0.130 0.925 0.650 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 2.740 4.100 3.000 ;
        RECT  1.715 2.525 1.975 3.000 ;
        RECT  0.925 2.740 1.715 3.000 ;
        RECT  0.665 2.525 0.925 3.000 ;
        RECT  0.000 2.740 0.665 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.815 0.565 3.975 2.395 ;
        RECT  3.645 0.565 3.815 0.825 ;
        RECT  3.715 1.795 3.815 2.395 ;
        RECT  0.930 2.185 3.715 2.345 ;
        RECT  2.745 0.475 2.905 2.005 ;
        RECT  2.675 0.475 2.745 0.825 ;
        RECT  1.465 0.475 2.675 0.635 ;
        RECT  2.495 1.270 2.565 1.530 ;
        RECT  2.335 0.815 2.495 1.915 ;
        RECT  2.115 0.815 2.335 0.975 ;
        RECT  2.185 1.755 2.335 1.915 ;
        RECT  1.365 0.380 1.465 0.980 ;
        RECT  1.365 1.745 1.465 2.005 ;
        RECT  1.205 0.380 1.365 2.005 ;
        RECT  0.930 1.225 1.010 1.485 ;
        RECT  0.770 0.830 0.930 2.345 ;
        RECT  0.385 0.830 0.770 0.990 ;
        RECT  0.385 2.185 0.770 2.345 ;
        RECT  0.125 0.385 0.385 0.990 ;
        RECT  0.125 1.825 0.385 2.425 ;
    END
END XNOR2X2MTH

MACRO XNOR2X4MTH
    CLASS CORE ;
    FOREIGN XNOR2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.530 1.785 5.615 2.385 ;
        RECT  5.350 0.345 5.530 2.385 ;
        RECT  5.245 0.345 5.350 0.880 ;
        RECT  4.490 0.345 5.245 0.525 ;
        RECT  4.490 1.785 4.595 2.045 ;
        RECT  4.310 0.345 4.490 2.210 ;
        RECT  4.200 0.345 4.310 1.170 ;
        RECT  3.585 2.030 4.310 2.210 ;
        RECT  3.405 0.715 3.585 2.210 ;
        RECT  3.205 0.715 3.405 0.875 ;
        RECT  3.315 1.710 3.405 1.970 ;
        END
        AntennaDiffArea 1.383 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.465 1.240 1.065 1.500 ;
        RECT  0.310 1.290 0.465 1.500 ;
        RECT  0.100 1.290 0.310 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.280 2.675 1.540 ;
        END
        AntennaGateArea 0.4862 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.455 -0.130 5.740 0.130 ;
        RECT  2.195 -0.130 2.455 0.250 ;
        RECT  1.405 -0.130 2.195 0.130 ;
        RECT  1.145 -0.130 1.405 0.650 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.980 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.515 2.740 5.740 3.000 ;
        RECT  2.255 2.510 2.515 3.000 ;
        RECT  1.435 2.740 2.255 3.000 ;
        RECT  1.175 2.510 1.435 3.000 ;
        RECT  0.385 2.740 1.175 3.000 ;
        RECT  0.125 1.805 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.895 0.705 5.055 2.560 ;
        RECT  4.735 0.705 4.895 0.965 ;
        RECT  3.045 2.400 4.895 2.560 ;
        RECT  3.925 1.690 4.085 1.850 ;
        RECT  3.765 0.375 3.925 1.850 ;
        RECT  2.995 0.375 3.765 0.535 ;
        RECT  3.025 1.230 3.225 1.490 ;
        RECT  3.025 1.720 3.065 1.980 ;
        RECT  2.885 2.170 3.045 2.560 ;
        RECT  2.865 0.770 3.025 1.980 ;
        RECT  2.835 0.375 2.995 0.590 ;
        RECT  1.470 2.170 2.885 2.330 ;
        RECT  2.695 0.770 2.865 0.930 ;
        RECT  2.805 1.720 2.865 1.980 ;
        RECT  1.925 0.430 2.835 0.590 ;
        RECT  1.915 0.430 1.925 1.990 ;
        RECT  1.765 0.375 1.915 1.990 ;
        RECT  1.655 0.375 1.765 0.975 ;
        RECT  1.470 1.225 1.585 1.485 ;
        RECT  1.310 0.830 1.470 2.330 ;
        RECT  0.895 0.830 1.310 0.990 ;
        RECT  0.895 2.170 1.310 2.330 ;
        RECT  0.635 0.390 0.895 0.990 ;
        RECT  0.635 1.805 0.895 2.405 ;
    END
END XNOR2X4MTH

MACRO XNOR2X8MTH
    CLASS CORE ;
    FOREIGN XNOR2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.660 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.425 1.810 10.535 2.410 ;
        RECT  10.165 0.310 10.425 2.410 ;
        RECT  9.475 0.310 10.165 0.525 ;
        RECT  9.475 1.945 9.515 2.205 ;
        RECT  9.215 0.310 9.475 2.205 ;
        RECT  9.145 0.310 9.215 0.825 ;
        RECT  8.505 0.310 9.145 0.525 ;
        RECT  8.505 1.085 8.550 2.220 ;
        RECT  8.165 0.310 8.505 2.220 ;
        RECT  7.475 2.030 8.165 2.220 ;
        RECT  7.215 0.715 7.475 2.220 ;
        RECT  7.100 0.715 7.215 0.875 ;
        RECT  6.460 2.030 7.215 2.220 ;
        RECT  6.300 0.715 6.460 2.220 ;
        RECT  6.080 0.715 6.300 0.875 ;
        RECT  6.195 1.805 6.300 2.220 ;
        END
        AntennaDiffArea 2.363 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.720 1.240 2.085 1.500 ;
        RECT  0.465 1.240 0.720 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.945 1.240 5.545 1.540 ;
        END
        AntennaGateArea 1.0062 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  4.835 -0.130 10.660 0.130 ;
        RECT  4.235 -0.130 4.835 0.250 ;
        RECT  3.445 -0.130 4.235 0.130 ;
        RECT  3.185 -0.130 3.445 0.675 ;
        RECT  2.425 -0.130 3.185 0.130 ;
        RECT  2.165 -0.130 2.425 0.635 ;
        RECT  1.405 -0.130 2.165 0.130 ;
        RECT  1.145 -0.130 1.405 0.650 ;
        RECT  0.385 -0.130 1.145 0.130 ;
        RECT  0.125 -0.130 0.385 0.965 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.345 2.740 10.660 3.000 ;
        RECT  4.405 2.620 5.345 3.000 ;
        RECT  3.535 2.740 4.405 3.000 ;
        RECT  3.275 2.425 3.535 3.000 ;
        RECT  2.455 2.740 3.275 3.000 ;
        RECT  2.195 2.425 2.455 3.000 ;
        RECT  1.405 2.740 2.195 3.000 ;
        RECT  1.145 2.180 1.405 3.000 ;
        RECT  0.385 2.740 1.145 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.815 0.705 9.975 2.560 ;
        RECT  9.655 0.705 9.815 0.965 ;
        RECT  9.005 2.400 9.815 2.560 ;
        RECT  8.955 1.815 9.005 2.560 ;
        RECT  8.795 0.705 8.955 2.560 ;
        RECT  8.685 0.705 8.795 0.965 ;
        RECT  8.745 1.815 8.795 2.560 ;
        RECT  5.965 2.400 8.745 2.560 ;
        RECT  7.825 1.690 7.985 1.850 ;
        RECT  7.665 0.375 7.825 1.850 ;
        RECT  6.800 0.375 7.665 0.535 ;
        RECT  6.800 1.690 6.965 1.850 ;
        RECT  6.640 0.375 6.800 1.850 ;
        RECT  5.905 0.375 6.640 0.535 ;
        RECT  5.945 1.230 6.120 1.490 ;
        RECT  5.805 2.085 5.965 2.560 ;
        RECT  5.900 1.230 5.945 1.905 ;
        RECT  5.745 0.375 5.905 0.590 ;
        RECT  5.740 0.770 5.900 1.905 ;
        RECT  3.495 2.085 5.805 2.245 ;
        RECT  4.425 0.430 5.745 0.590 ;
        RECT  4.605 0.770 5.740 0.930 ;
        RECT  4.725 1.745 5.740 1.905 ;
        RECT  4.265 0.430 4.425 1.895 ;
        RECT  3.955 0.860 4.265 1.020 ;
        RECT  3.815 1.735 4.265 1.895 ;
        RECT  3.495 1.225 4.020 1.485 ;
        RECT  3.695 0.385 3.955 1.020 ;
        RECT  2.935 0.860 3.695 1.020 ;
        RECT  3.335 1.225 3.495 2.245 ;
        RECT  3.080 1.225 3.335 1.485 ;
        RECT  2.460 2.085 3.335 2.245 ;
        RECT  2.835 1.735 2.995 1.895 ;
        RECT  2.835 0.420 2.935 1.020 ;
        RECT  2.675 0.420 2.835 1.895 ;
        RECT  2.300 0.830 2.460 2.245 ;
        RECT  1.915 0.830 2.300 0.990 ;
        RECT  1.915 1.840 2.300 2.000 ;
        RECT  1.655 0.390 1.915 0.990 ;
        RECT  1.655 1.840 1.915 2.455 ;
        RECT  0.895 0.830 1.655 0.990 ;
        RECT  0.895 1.840 1.655 2.000 ;
        RECT  0.635 0.380 0.895 0.990 ;
        RECT  0.635 1.840 0.895 2.460 ;
    END
END XNOR2X8MTH

MACRO XNOR2XLMTH
    CLASS CORE ;
    FOREIGN XNOR2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.495 1.290 3.590 1.580 ;
        RECT  3.235 0.765 3.495 1.945 ;
        RECT  3.175 0.765 3.235 1.025 ;
        END
        AntennaDiffArea 0.238 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.505 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.645 1.215 2.065 1.580 ;
        END
        AntennaGateArea 0.1066 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.680 -0.130 4.100 0.130 ;
        RECT  0.740 -0.130 1.680 0.295 ;
        RECT  0.000 -0.130 0.740 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.745 2.740 4.100 3.000 ;
        RECT  0.805 2.465 1.745 3.000 ;
        RECT  0.000 2.740 0.805 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.815 0.335 3.975 2.515 ;
        RECT  3.715 0.335 3.815 0.595 ;
        RECT  3.715 2.125 3.815 2.515 ;
        RECT  0.930 2.125 3.715 2.285 ;
        RECT  2.785 0.475 2.945 1.945 ;
        RECT  2.605 0.475 2.785 1.025 ;
        RECT  2.665 1.685 2.785 1.945 ;
        RECT  1.415 0.475 2.605 0.635 ;
        RECT  2.415 1.255 2.575 1.515 ;
        RECT  2.255 0.815 2.415 1.920 ;
        RECT  2.095 0.815 2.255 0.975 ;
        RECT  2.155 1.760 2.255 1.920 ;
        RECT  1.255 0.475 1.415 1.945 ;
        RECT  1.165 0.765 1.255 1.025 ;
        RECT  1.135 1.685 1.255 1.945 ;
        RECT  0.930 1.225 1.055 1.485 ;
        RECT  0.770 0.865 0.930 2.285 ;
        RECT  0.385 0.865 0.770 1.025 ;
        RECT  0.155 1.760 0.770 1.920 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END XNOR2XLMTH

MACRO XNOR3X1MTH
    CLASS CORE ;
    FOREIGN XNOR3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.050 0.755 8.100 1.580 ;
        RECT  8.050 2.170 8.075 2.330 ;
        RECT  7.890 0.755 8.050 2.330 ;
        RECT  7.865 0.755 7.890 1.015 ;
        RECT  7.815 2.170 7.890 2.330 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.635 1.700 7.690 1.990 ;
        RECT  7.475 1.700 7.635 2.405 ;
        RECT  7.095 2.245 7.475 2.405 ;
        RECT  6.835 2.245 7.095 2.445 ;
        END
        AntennaGateArea 0.1976 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 1.020 4.820 1.740 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.450 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.910 -0.130 8.200 0.130 ;
        RECT  7.310 -0.130 7.910 0.250 ;
        RECT  4.830 -0.130 7.310 0.130 ;
        RECT  4.610 -0.130 4.830 0.840 ;
        RECT  2.810 -0.130 4.610 0.130 ;
        RECT  2.650 -0.130 2.810 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 2.740 8.200 3.000 ;
        RECT  7.275 2.585 7.535 3.000 ;
        RECT  4.820 2.740 7.275 3.000 ;
        RECT  4.595 2.265 4.820 3.000 ;
        RECT  2.545 2.740 4.595 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.685 1.260 7.710 1.520 ;
        RECT  7.525 0.430 7.685 1.520 ;
        RECT  7.095 0.430 7.525 0.590 ;
        RECT  6.935 0.310 7.095 0.590 ;
        RECT  6.860 1.905 7.080 2.065 ;
        RECT  6.860 0.815 7.000 0.975 ;
        RECT  5.930 0.310 6.935 0.470 ;
        RECT  6.700 0.815 6.860 2.065 ;
        RECT  6.650 1.145 6.700 1.405 ;
        RECT  6.440 1.980 6.520 2.240 ;
        RECT  6.440 0.785 6.490 1.045 ;
        RECT  6.280 0.785 6.440 2.560 ;
        RECT  6.230 0.785 6.280 1.045 ;
        RECT  5.160 2.400 6.280 2.560 ;
        RECT  5.930 1.860 6.060 2.120 ;
        RECT  5.770 0.310 5.930 2.120 ;
        RECT  5.430 0.655 5.590 2.135 ;
        RECT  5.210 0.655 5.430 0.915 ;
        RECT  5.340 1.875 5.430 2.135 ;
        RECT  5.160 1.315 5.250 1.575 ;
        RECT  5.000 1.315 5.160 2.560 ;
        RECT  4.415 1.925 5.000 2.085 ;
        RECT  4.270 0.310 4.430 1.745 ;
        RECT  4.255 1.925 4.415 2.560 ;
        RECT  3.430 0.310 4.270 0.470 ;
        RECT  4.075 1.585 4.270 1.745 ;
        RECT  2.885 2.400 4.255 2.560 ;
        RECT  3.930 0.655 4.090 1.385 ;
        RECT  3.915 1.585 4.075 2.220 ;
        RECT  3.735 1.225 3.930 1.385 ;
        RECT  3.225 2.060 3.915 2.220 ;
        RECT  2.470 0.885 3.750 1.045 ;
        RECT  3.575 1.225 3.735 1.880 ;
        RECT  1.875 1.225 3.575 1.385 ;
        RECT  3.170 0.310 3.430 0.675 ;
        RECT  3.065 1.565 3.225 2.220 ;
        RECT  1.865 1.565 3.065 1.725 ;
        RECT  2.725 1.905 2.885 2.560 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.895 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.675 2.130 0.935 ;
        RECT  1.405 2.320 2.045 2.480 ;
        RECT  1.695 0.775 1.970 0.935 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.355 1.875 1.405 2.480 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  1.145 1.875 1.195 2.480 ;
        RECT  0.845 0.310 0.895 0.720 ;
        RECT  0.845 1.810 0.895 2.410 ;
        RECT  0.685 0.310 0.845 2.410 ;
        RECT  0.635 0.460 0.685 0.720 ;
        RECT  0.635 1.810 0.685 2.410 ;
    END
END XNOR3X1MTH

MACRO XNOR3X2MTH
    CLASS CORE ;
    FOREIGN XNOR3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.940 0.415 8.100 2.065 ;
        RECT  7.865 0.415 7.940 1.170 ;
        RECT  7.865 1.805 7.940 2.065 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.480 2.110 7.690 2.410 ;
        RECT  6.700 2.250 7.480 2.410 ;
        END
        AntennaGateArea 0.2444 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.075 4.820 1.745 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.450 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 -0.130 8.200 0.130 ;
        RECT  7.275 -0.130 7.535 0.250 ;
        RECT  4.840 -0.130 7.275 0.130 ;
        RECT  4.580 -0.130 4.840 0.835 ;
        RECT  2.870 -0.130 4.580 0.130 ;
        RECT  2.650 -0.130 2.870 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 2.740 8.200 3.000 ;
        RECT  7.275 2.595 7.535 3.000 ;
        RECT  4.820 2.740 7.275 3.000 ;
        RECT  4.595 2.265 4.820 3.000 ;
        RECT  2.545 2.740 4.595 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.685 1.265 7.710 1.525 ;
        RECT  7.525 0.430 7.685 1.525 ;
        RECT  5.900 0.430 7.525 0.590 ;
        RECT  6.860 1.875 7.080 2.035 ;
        RECT  6.860 0.815 6.970 0.975 ;
        RECT  6.700 0.815 6.860 2.035 ;
        RECT  6.620 1.165 6.700 1.425 ;
        RECT  6.400 1.835 6.520 2.435 ;
        RECT  6.400 0.840 6.460 1.000 ;
        RECT  6.240 0.840 6.400 2.560 ;
        RECT  6.200 0.840 6.240 1.000 ;
        RECT  5.160 2.400 6.240 2.560 ;
        RECT  5.900 1.855 6.060 2.115 ;
        RECT  5.740 0.430 5.900 2.115 ;
        RECT  5.400 0.630 5.560 2.140 ;
        RECT  5.230 0.630 5.400 0.890 ;
        RECT  5.340 1.880 5.400 2.140 ;
        RECT  5.160 1.265 5.220 1.525 ;
        RECT  5.000 1.265 5.160 2.560 ;
        RECT  4.415 1.925 5.000 2.085 ;
        RECT  4.255 1.925 4.415 2.560 ;
        RECT  4.240 0.310 4.400 1.745 ;
        RECT  2.885 2.400 4.255 2.560 ;
        RECT  3.435 0.310 4.240 0.470 ;
        RECT  4.075 1.585 4.240 1.745 ;
        RECT  3.915 1.585 4.075 2.220 ;
        RECT  3.900 0.665 4.060 1.385 ;
        RECT  3.225 2.060 3.915 2.220 ;
        RECT  3.735 1.225 3.900 1.385 ;
        RECT  3.575 1.225 3.735 1.880 ;
        RECT  2.470 0.885 3.720 1.045 ;
        RECT  1.875 1.225 3.575 1.385 ;
        RECT  3.175 0.310 3.435 0.675 ;
        RECT  3.065 1.565 3.225 2.220 ;
        RECT  1.865 1.565 3.065 1.725 ;
        RECT  2.725 1.905 2.885 2.560 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.845 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.675 2.130 0.935 ;
        RECT  1.355 2.320 2.045 2.480 ;
        RECT  1.695 0.775 1.970 0.935 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  0.685 0.310 0.845 2.415 ;
    END
END XNOR3X2MTH

MACRO XNOR3X4MTH
    CLASS CORE ;
    FOREIGN XNOR3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.685 0.415 8.865 2.410 ;
        RECT  8.535 0.415 8.685 1.015 ;
        RECT  8.535 1.700 8.685 2.410 ;
        RECT  8.300 1.700 8.535 1.990 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.890 2.110 8.100 2.405 ;
        RECT  7.250 2.245 7.890 2.405 ;
        END
        AntennaGateArea 0.2444 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.545 1.120 4.820 1.580 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.500 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 -0.130 9.430 0.130 ;
        RECT  9.045 -0.130 9.305 1.015 ;
        RECT  8.255 -0.130 9.045 0.130 ;
        RECT  7.995 -0.130 8.255 0.250 ;
        RECT  5.590 -0.130 7.995 0.130 ;
        RECT  5.340 -0.130 5.590 0.745 ;
        RECT  2.825 -0.130 5.340 0.130 ;
        RECT  2.665 -0.130 2.825 0.705 ;
        RECT  0.385 -0.130 2.665 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 2.740 9.430 3.000 ;
        RECT  9.045 1.830 9.305 3.000 ;
        RECT  8.255 2.740 9.045 3.000 ;
        RECT  7.995 2.595 8.255 3.000 ;
        RECT  5.560 2.740 7.995 3.000 ;
        RECT  5.300 2.605 5.560 3.000 ;
        RECT  2.580 2.740 5.300 3.000 ;
        RECT  2.420 2.245 2.580 3.000 ;
        RECT  0.385 2.740 2.420 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.355 1.235 8.505 1.495 ;
        RECT  8.195 0.430 8.355 1.495 ;
        RECT  6.560 0.430 8.195 0.590 ;
        RECT  7.530 1.875 7.660 2.035 ;
        RECT  7.530 0.815 7.630 0.975 ;
        RECT  7.370 0.815 7.530 2.035 ;
        RECT  7.250 1.245 7.370 1.505 ;
        RECT  7.070 0.840 7.120 1.000 ;
        RECT  6.910 0.840 7.070 2.425 ;
        RECT  6.860 0.840 6.910 1.000 ;
        RECT  5.500 2.265 6.910 2.425 ;
        RECT  6.400 0.430 6.560 2.085 ;
        RECT  6.020 0.630 6.180 2.085 ;
        RECT  5.890 0.630 6.020 1.085 ;
        RECT  5.890 1.825 6.020 2.085 ;
        RECT  5.160 0.925 5.890 1.085 ;
        RECT  5.500 1.265 5.840 1.525 ;
        RECT  5.340 1.265 5.500 2.425 ;
        RECT  4.530 2.265 5.340 2.425 ;
        RECT  5.000 0.615 5.160 2.045 ;
        RECT  4.820 0.615 5.000 0.875 ;
        RECT  4.760 1.885 5.000 2.045 ;
        RECT  4.370 2.265 4.530 2.560 ;
        RECT  2.920 2.400 4.370 2.560 ;
        RECT  4.205 0.310 4.365 1.745 ;
        RECT  3.445 0.310 4.205 0.470 ;
        RECT  4.190 1.585 4.205 1.745 ;
        RECT  4.030 1.585 4.190 2.220 ;
        RECT  3.340 2.060 4.030 2.220 ;
        RECT  3.865 0.650 4.025 1.385 ;
        RECT  3.850 1.225 3.865 1.385 ;
        RECT  3.690 1.225 3.850 1.880 ;
        RECT  1.875 1.225 3.690 1.385 ;
        RECT  2.485 0.885 3.685 1.045 ;
        RECT  3.185 0.310 3.445 0.675 ;
        RECT  3.180 1.565 3.340 2.220 ;
        RECT  1.900 1.565 3.180 1.725 ;
        RECT  2.760 1.905 2.920 2.560 ;
        RECT  2.240 1.905 2.760 2.065 ;
        RECT  2.325 0.310 2.485 1.045 ;
        RECT  0.895 0.310 2.325 0.470 ;
        RECT  2.080 1.905 2.240 2.480 ;
        RECT  1.985 0.675 2.145 0.935 ;
        RECT  1.355 2.320 2.080 2.480 ;
        RECT  1.695 0.775 1.985 0.935 ;
        RECT  1.740 1.565 1.900 2.140 ;
        RECT  1.695 1.565 1.740 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  0.845 0.310 0.895 0.815 ;
        RECT  0.685 0.310 0.845 2.410 ;
        RECT  0.635 0.310 0.685 0.815 ;
    END
END XNOR3X4MTH

MACRO XNOR3X8MTH
    CLASS CORE ;
    FOREIGN XNOR3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.480 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.540 0.415 10.890 2.450 ;
        RECT  10.105 0.745 10.540 2.025 ;
        RECT  9.850 0.745 10.105 1.055 ;
        RECT  9.870 1.675 10.105 2.025 ;
        RECT  9.520 1.675 9.870 2.450 ;
        RECT  9.540 0.415 9.850 1.055 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  9.075 1.700 9.330 1.990 ;
        RECT  8.915 1.700 9.075 2.410 ;
        RECT  8.630 2.250 8.915 2.410 ;
        END
        AntennaGateArea 0.2444 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.120 5.030 1.580 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.500 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.345 -0.130 11.480 0.130 ;
        RECT  11.105 -0.130 11.345 0.990 ;
        RECT  10.335 -0.130 11.105 0.130 ;
        RECT  10.075 -0.130 10.335 0.565 ;
        RECT  9.285 -0.130 10.075 0.130 ;
        RECT  9.025 -0.130 9.285 0.295 ;
        RECT  6.650 -0.130 9.025 0.130 ;
        RECT  6.390 -0.130 6.650 0.565 ;
        RECT  5.630 -0.130 6.390 0.130 ;
        RECT  5.370 -0.130 5.630 0.565 ;
        RECT  2.810 -0.130 5.370 0.130 ;
        RECT  2.650 -0.130 2.810 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  11.345 2.740 11.480 3.000 ;
        RECT  11.105 1.825 11.345 3.000 ;
        RECT  10.335 2.740 11.105 3.000 ;
        RECT  10.075 2.205 10.335 3.000 ;
        RECT  9.285 2.740 10.075 3.000 ;
        RECT  9.025 2.620 9.285 3.000 ;
        RECT  6.630 2.740 9.025 3.000 ;
        RECT  6.370 2.570 6.630 3.000 ;
        RECT  5.510 2.740 6.370 3.000 ;
        RECT  5.250 2.570 5.510 3.000 ;
        RECT  2.545 2.740 5.250 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  9.270 1.235 9.925 1.495 ;
        RECT  9.110 0.475 9.270 1.495 ;
        RECT  7.620 0.475 9.110 0.635 ;
        RECT  8.430 0.815 8.720 2.035 ;
        RECT  8.215 1.335 8.430 1.595 ;
        RECT  8.035 1.835 8.210 2.435 ;
        RECT  8.035 0.845 8.180 1.105 ;
        RECT  7.875 0.845 8.035 2.435 ;
        RECT  7.215 2.275 7.875 2.435 ;
        RECT  7.620 1.825 7.650 2.085 ;
        RECT  7.460 0.475 7.620 2.085 ;
        RECT  7.120 0.645 7.280 2.035 ;
        RECT  7.055 2.230 7.215 2.435 ;
        RECT  6.900 0.645 7.120 0.905 ;
        RECT  6.925 1.775 7.120 2.035 ;
        RECT  6.660 2.230 7.055 2.390 ;
        RECT  6.140 0.745 6.900 0.905 ;
        RECT  6.500 1.265 6.660 2.390 ;
        RECT  5.700 1.265 6.500 1.525 ;
        RECT  4.415 2.230 6.500 2.390 ;
        RECT  5.880 0.575 6.140 0.905 ;
        RECT  5.430 1.885 6.090 2.045 ;
        RECT  5.430 0.745 5.880 0.905 ;
        RECT  5.270 0.745 5.430 2.045 ;
        RECT  5.120 0.745 5.270 0.905 ;
        RECT  4.670 1.885 5.270 2.045 ;
        RECT  4.860 0.540 5.120 0.905 ;
        RECT  4.255 2.230 4.415 2.560 ;
        RECT  4.240 0.310 4.400 1.745 ;
        RECT  2.885 2.400 4.255 2.560 ;
        RECT  3.430 0.310 4.240 0.470 ;
        RECT  4.075 1.585 4.240 1.745 ;
        RECT  3.915 1.585 4.075 2.220 ;
        RECT  3.900 0.650 4.060 1.385 ;
        RECT  3.225 2.060 3.915 2.220 ;
        RECT  3.735 1.225 3.900 1.385 ;
        RECT  3.575 1.225 3.735 1.880 ;
        RECT  2.470 0.885 3.720 1.045 ;
        RECT  1.875 1.225 3.575 1.385 ;
        RECT  3.170 0.310 3.430 0.675 ;
        RECT  3.065 1.565 3.225 2.220 ;
        RECT  1.865 1.565 3.065 1.725 ;
        RECT  2.725 1.905 2.885 2.560 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.845 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.675 2.130 0.935 ;
        RECT  1.355 2.320 2.045 2.480 ;
        RECT  1.695 0.775 1.970 0.935 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  0.845 1.810 0.895 2.410 ;
        RECT  0.685 0.310 0.845 2.410 ;
        RECT  0.635 1.810 0.685 2.410 ;
    END
END XNOR3X8MTH

MACRO XNOR3XLMTH
    CLASS CORE ;
    FOREIGN XNOR3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.890 0.765 8.100 1.930 ;
        RECT  7.865 0.765 7.890 1.025 ;
        RECT  7.815 1.770 7.890 1.930 ;
        END
        AntennaDiffArea 0.225 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.480 2.110 7.690 2.400 ;
        RECT  6.700 2.165 7.480 2.400 ;
        END
        AntennaGateArea 0.169 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.610 1.020 4.820 1.740 ;
        END
        AntennaGateArea 0.1794 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.500 1.580 ;
        END
        AntennaGateArea 0.1378 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.910 -0.130 8.200 0.130 ;
        RECT  7.310 -0.130 7.910 0.295 ;
        RECT  4.830 -0.130 7.310 0.130 ;
        RECT  4.610 -0.130 4.830 0.840 ;
        RECT  2.810 -0.130 4.610 0.130 ;
        RECT  2.650 -0.130 2.810 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.835 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.990 2.740 8.200 3.000 ;
        RECT  7.390 2.585 7.990 3.000 ;
        RECT  4.820 2.740 7.390 3.000 ;
        RECT  4.595 2.265 4.820 3.000 ;
        RECT  2.545 2.740 4.595 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.985 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.685 1.260 7.710 1.520 ;
        RECT  7.525 0.475 7.685 1.520 ;
        RECT  7.095 0.475 7.525 0.635 ;
        RECT  6.935 0.310 7.095 0.635 ;
        RECT  6.860 1.805 7.080 1.965 ;
        RECT  6.860 0.815 7.000 0.975 ;
        RECT  5.930 0.310 6.935 0.470 ;
        RECT  6.700 0.815 6.860 1.965 ;
        RECT  6.650 1.195 6.700 1.455 ;
        RECT  6.440 1.980 6.520 2.240 ;
        RECT  6.440 0.785 6.490 1.045 ;
        RECT  6.280 0.785 6.440 2.560 ;
        RECT  6.230 0.785 6.280 1.045 ;
        RECT  5.160 2.400 6.280 2.560 ;
        RECT  5.930 1.855 6.060 2.115 ;
        RECT  5.770 0.310 5.930 2.115 ;
        RECT  5.430 0.655 5.590 2.115 ;
        RECT  5.210 0.655 5.430 0.915 ;
        RECT  5.340 1.855 5.430 2.115 ;
        RECT  5.160 1.315 5.250 1.575 ;
        RECT  5.000 1.315 5.160 2.560 ;
        RECT  4.415 1.925 5.000 2.085 ;
        RECT  4.270 0.310 4.430 1.745 ;
        RECT  4.255 1.925 4.415 2.560 ;
        RECT  3.430 0.310 4.270 0.470 ;
        RECT  4.075 1.585 4.270 1.745 ;
        RECT  2.885 2.400 4.255 2.560 ;
        RECT  3.930 0.655 4.090 1.385 ;
        RECT  3.915 1.585 4.075 2.220 ;
        RECT  3.735 1.225 3.930 1.385 ;
        RECT  3.225 2.060 3.915 2.220 ;
        RECT  2.470 0.885 3.750 1.045 ;
        RECT  3.575 1.225 3.735 1.880 ;
        RECT  1.875 1.225 3.575 1.385 ;
        RECT  3.170 0.310 3.430 0.675 ;
        RECT  3.065 1.565 3.225 2.220 ;
        RECT  1.865 1.565 3.065 1.725 ;
        RECT  2.725 1.905 2.885 2.560 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.845 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.675 2.130 0.935 ;
        RECT  1.355 2.320 2.045 2.480 ;
        RECT  1.695 0.775 1.970 0.935 ;
        RECT  1.705 1.565 1.865 2.115 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  0.685 0.310 0.845 2.245 ;
    END
END XNOR3XLMTH

MACRO XOR2X1MTH
    CLASS CORE ;
    FOREIGN XOR2X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.465 1.290 3.590 1.580 ;
        RECT  3.355 1.290 3.465 1.945 ;
        RECT  3.305 0.765 3.355 1.945 ;
        RECT  3.195 0.765 3.305 1.450 ;
        RECT  3.205 1.685 3.305 1.945 ;
        RECT  3.095 0.765 3.195 1.025 ;
        END
        AntennaDiffArea 0.258 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.200 0.555 1.580 ;
        END
        AntennaGateArea 0.1274 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.550 1.215 1.950 1.830 ;
        END
        AntennaGateArea 0.1417 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  3.890 -0.130 4.100 0.130 ;
        RECT  2.950 -0.130 3.890 0.280 ;
        RECT  2.580 -0.130 2.950 0.130 ;
        RECT  1.980 -0.130 2.580 0.280 ;
        RECT  1.605 -0.130 1.980 0.130 ;
        RECT  0.665 -0.130 1.605 0.280 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.865 2.740 4.100 3.000 ;
        RECT  0.925 2.555 1.865 3.000 ;
        RECT  0.540 2.740 0.925 3.000 ;
        RECT  0.280 2.555 0.540 3.000 ;
        RECT  0.000 2.740 0.280 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.930 1.765 3.975 2.025 ;
        RECT  3.770 0.765 3.930 2.285 ;
        RECT  3.605 0.765 3.770 1.025 ;
        RECT  3.715 1.765 3.770 2.285 ;
        RECT  1.325 2.125 3.715 2.285 ;
        RECT  2.910 1.685 2.955 1.945 ;
        RECT  2.750 0.475 2.910 1.945 ;
        RECT  2.585 0.475 2.750 1.025 ;
        RECT  2.695 1.685 2.750 1.945 ;
        RECT  0.935 0.475 2.585 0.635 ;
        RECT  2.405 1.245 2.570 1.505 ;
        RECT  2.405 1.760 2.445 1.920 ;
        RECT  2.245 0.815 2.405 1.920 ;
        RECT  2.075 0.815 2.245 0.975 ;
        RECT  2.185 1.760 2.245 1.920 ;
        RECT  1.325 0.815 1.375 0.975 ;
        RECT  1.165 0.815 1.325 2.285 ;
        RECT  1.115 0.815 1.165 0.975 ;
        RECT  0.935 1.225 0.985 1.485 ;
        RECT  0.775 0.475 0.935 1.920 ;
        RECT  0.385 0.830 0.775 0.990 ;
        RECT  0.385 1.760 0.775 1.920 ;
        RECT  0.125 0.730 0.385 0.990 ;
        RECT  0.125 1.760 0.385 2.020 ;
    END
END XOR2X1MTH

MACRO XOR2X2MTH
    CLASS CORE ;
    FOREIGN XOR2X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.365 1.290 3.590 1.580 ;
        RECT  3.365 1.865 3.465 2.025 ;
        RECT  3.365 0.560 3.395 0.820 ;
        RECT  3.205 0.560 3.365 2.025 ;
        RECT  3.135 0.560 3.205 0.820 ;
        END
        AntennaDiffArea 0.499 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.290 0.555 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.985 1.155 2.090 1.525 ;
        RECT  1.645 1.155 1.985 1.580 ;
        END
        AntennaGateArea 0.2522 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.975 -0.130 4.100 0.130 ;
        RECT  1.715 -0.130 1.975 0.290 ;
        RECT  0.925 -0.130 1.715 0.130 ;
        RECT  0.665 -0.130 0.925 0.250 ;
        RECT  0.000 -0.130 0.665 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.915 2.740 4.100 3.000 ;
        RECT  1.655 2.545 1.915 3.000 ;
        RECT  0.895 2.740 1.655 3.000 ;
        RECT  0.635 2.170 0.895 3.000 ;
        RECT  0.000 2.740 0.635 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.815 0.560 3.975 2.365 ;
        RECT  3.645 0.560 3.815 0.820 ;
        RECT  3.715 1.815 3.815 2.365 ;
        RECT  1.465 2.205 3.715 2.365 ;
        RECT  2.795 0.475 2.955 2.025 ;
        RECT  2.675 0.475 2.795 0.820 ;
        RECT  2.695 1.765 2.795 2.025 ;
        RECT  0.965 0.475 2.675 0.635 ;
        RECT  2.465 1.270 2.615 1.530 ;
        RECT  2.305 0.815 2.465 1.965 ;
        RECT  2.115 0.815 2.305 0.975 ;
        RECT  2.185 1.705 2.305 1.965 ;
        RECT  1.405 0.815 1.465 2.365 ;
        RECT  1.305 0.815 1.405 2.485 ;
        RECT  1.205 0.815 1.305 0.975 ;
        RECT  1.145 1.885 1.305 2.485 ;
        RECT  0.965 1.240 1.125 1.500 ;
        RECT  0.805 0.475 0.965 1.930 ;
        RECT  0.385 0.830 0.805 0.990 ;
        RECT  0.385 1.770 0.805 1.930 ;
        RECT  0.125 0.390 0.385 0.990 ;
        RECT  0.125 1.770 0.385 2.370 ;
    END
END XOR2X2MTH

MACRO XOR2X3MTH
    CLASS CORE ;
    FOREIGN XOR2X3MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.495 1.820 5.605 2.080 ;
        RECT  5.335 0.355 5.495 2.080 ;
        RECT  5.235 0.355 5.335 0.880 ;
        RECT  4.475 0.355 5.235 0.515 ;
        RECT  4.425 0.355 4.475 0.885 ;
        RECT  4.425 1.820 4.475 2.080 ;
        RECT  4.200 0.355 4.425 2.205 ;
        RECT  3.475 2.045 4.200 2.205 ;
        RECT  3.315 0.715 3.475 2.205 ;
        RECT  3.195 0.715 3.315 0.875 ;
        RECT  3.245 1.710 3.315 1.970 ;
        END
        AntennaDiffArea 1.162 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.290 1.095 1.450 ;
        RECT  0.100 1.290 0.310 1.580 ;
        END
        AntennaGateArea 0.312 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.110 1.295 2.605 1.555 ;
        END
        AntennaGateArea 0.377 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 -0.130 5.740 0.130 ;
        RECT  2.285 -0.130 2.545 0.250 ;
        RECT  1.465 -0.130 2.285 0.130 ;
        RECT  1.205 -0.130 1.465 0.250 ;
        RECT  0.385 -0.130 1.205 0.130 ;
        RECT  0.125 -0.130 0.385 0.990 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.545 2.740 5.740 3.000 ;
        RECT  2.285 2.510 2.545 3.000 ;
        RECT  1.465 2.740 2.285 3.000 ;
        RECT  1.205 2.040 1.465 3.000 ;
        RECT  0.385 2.740 1.205 3.000 ;
        RECT  0.125 1.770 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  4.995 1.820 5.095 2.080 ;
        RECT  4.835 0.705 4.995 2.545 ;
        RECT  4.725 0.705 4.835 0.965 ;
        RECT  3.045 2.385 4.835 2.545 ;
        RECT  3.865 0.625 3.965 0.885 ;
        RECT  3.865 1.705 3.965 1.865 ;
        RECT  3.705 0.375 3.865 1.865 ;
        RECT  2.995 0.375 3.705 0.535 ;
        RECT  2.970 1.230 3.135 1.490 ;
        RECT  2.885 2.170 3.045 2.545 ;
        RECT  2.835 0.375 2.995 0.590 ;
        RECT  2.810 0.770 2.970 1.905 ;
        RECT  1.955 2.170 2.885 2.330 ;
        RECT  1.470 0.430 2.835 0.590 ;
        RECT  2.685 0.770 2.810 0.930 ;
        RECT  2.685 1.745 2.810 1.905 ;
        RECT  1.930 0.815 2.005 0.975 ;
        RECT  1.930 1.700 1.955 2.330 ;
        RECT  1.770 0.815 1.930 2.330 ;
        RECT  1.745 0.815 1.770 0.975 ;
        RECT  1.470 1.225 1.590 1.485 ;
        RECT  1.310 0.430 1.470 1.860 ;
        RECT  0.925 0.745 1.310 0.905 ;
        RECT  0.925 1.700 1.310 1.860 ;
        RECT  0.665 0.645 0.925 0.905 ;
        RECT  0.665 1.700 0.925 2.300 ;
    END
END XOR2X3MTH

MACRO XOR2X4MTH
    CLASS CORE ;
    FOREIGN XOR2X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.740 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.505 1.745 5.615 2.345 ;
        RECT  5.345 0.370 5.505 2.345 ;
        RECT  5.245 0.370 5.345 0.835 ;
        RECT  4.495 0.370 5.245 0.530 ;
        RECT  4.495 1.815 4.595 2.205 ;
        RECT  4.335 0.370 4.495 2.205 ;
        RECT  4.225 0.370 4.335 0.835 ;
        RECT  4.160 1.330 4.335 1.540 ;
        RECT  3.525 2.045 4.335 2.205 ;
        RECT  3.365 0.770 3.525 2.205 ;
        RECT  3.205 0.770 3.365 0.930 ;
        END
        AntennaDiffArea 1.39 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.310 1.240 1.065 1.500 ;
        RECT  0.100 1.240 0.310 1.580 ;
        END
        AntennaGateArea 0.4108 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  2.150 1.245 2.685 1.580 ;
        END
        AntennaGateArea 0.4862 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.525 -0.130 5.740 0.130 ;
        RECT  2.265 -0.130 2.525 0.250 ;
        RECT  1.445 -0.130 2.265 0.130 ;
        RECT  1.185 -0.130 1.445 0.250 ;
        RECT  0.385 -0.130 1.185 0.130 ;
        RECT  0.125 -0.130 0.385 0.990 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  2.525 2.740 5.740 3.000 ;
        RECT  2.265 2.540 2.525 3.000 ;
        RECT  1.440 2.740 2.265 3.000 ;
        RECT  1.180 2.070 1.440 3.000 ;
        RECT  0.385 2.740 1.180 3.000 ;
        RECT  0.125 1.905 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  5.005 1.745 5.105 2.345 ;
        RECT  4.845 0.720 5.005 2.545 ;
        RECT  4.735 0.720 4.845 0.980 ;
        RECT  3.045 2.385 4.845 2.545 ;
        RECT  3.980 1.705 4.085 1.865 ;
        RECT  3.820 0.375 3.980 1.865 ;
        RECT  3.715 0.375 3.820 0.835 ;
        RECT  3.165 0.375 3.715 0.535 ;
        RECT  3.065 1.230 3.185 1.490 ;
        RECT  3.005 0.375 3.165 0.590 ;
        RECT  3.025 1.230 3.065 2.005 ;
        RECT  2.885 2.200 3.045 2.545 ;
        RECT  2.865 0.770 3.025 2.005 ;
        RECT  1.545 0.430 3.005 0.590 ;
        RECT  1.935 2.200 2.885 2.360 ;
        RECT  2.695 0.770 2.865 0.930 ;
        RECT  2.805 1.745 2.865 2.005 ;
        RECT  1.935 0.770 1.985 0.930 ;
        RECT  1.775 0.770 1.935 2.360 ;
        RECT  1.725 0.770 1.775 0.930 ;
        RECT  1.545 1.225 1.595 1.485 ;
        RECT  1.385 0.430 1.545 1.890 ;
        RECT  0.895 0.830 1.385 0.990 ;
        RECT  0.895 1.730 1.385 1.890 ;
        RECT  0.635 0.390 0.895 0.990 ;
        RECT  0.635 1.730 0.895 2.400 ;
    END
END XOR2X4MTH

MACRO XOR2X8MTH
    CLASS CORE ;
    FOREIGN XOR2X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.810 1.810 10.945 2.410 ;
        RECT  10.600 0.310 10.810 2.410 ;
        RECT  9.790 0.310 10.600 0.520 ;
        RECT  9.790 1.960 9.925 2.220 ;
        RECT  9.580 0.310 9.790 2.220 ;
        RECT  8.915 0.310 9.580 0.520 ;
        RECT  8.915 1.085 8.960 2.220 ;
        RECT  8.575 0.310 8.915 2.220 ;
        RECT  7.830 2.030 8.575 2.220 ;
        RECT  7.670 0.755 7.830 2.220 ;
        RECT  7.510 0.755 7.670 0.915 ;
        RECT  6.870 2.030 7.670 2.220 ;
        RECT  6.680 0.715 6.870 2.220 ;
        RECT  6.490 0.715 6.680 0.930 ;
        RECT  6.605 1.710 6.680 2.220 ;
        END
        AntennaDiffArea 2.365 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.130 1.240 2.130 1.500 ;
        RECT  0.510 1.240 1.130 1.580 ;
        END
        AntennaGateArea 0.8216 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.385 1.240 5.970 1.540 ;
        END
        AntennaGateArea 1.0062 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.700 -0.130 11.070 0.130 ;
        RECT  5.440 -0.130 5.700 0.250 ;
        RECT  4.720 -0.130 5.440 0.130 ;
        RECT  4.460 -0.130 4.720 0.250 ;
        RECT  3.640 -0.130 4.460 0.130 ;
        RECT  3.380 -0.130 3.640 0.290 ;
        RECT  2.560 -0.130 3.380 0.130 ;
        RECT  2.300 -0.130 2.560 0.290 ;
        RECT  1.480 -0.130 2.300 0.130 ;
        RECT  1.220 -0.130 1.480 0.650 ;
        RECT  0.400 -0.130 1.220 0.130 ;
        RECT  0.140 -0.130 0.400 1.025 ;
        RECT  0.000 -0.130 0.140 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  5.760 2.740 11.070 3.000 ;
        RECT  5.600 2.425 5.760 3.000 ;
        RECT  5.400 2.740 5.600 3.000 ;
        RECT  4.460 2.620 5.400 3.000 ;
        RECT  3.640 2.740 4.460 3.000 ;
        RECT  3.380 2.080 3.640 3.000 ;
        RECT  2.560 2.740 3.380 3.000 ;
        RECT  2.300 2.100 2.560 3.000 ;
        RECT  1.480 2.740 2.300 3.000 ;
        RECT  1.220 2.180 1.480 3.000 ;
        RECT  0.400 2.740 1.220 3.000 ;
        RECT  0.140 1.725 0.400 3.000 ;
        RECT  0.000 2.740 0.140 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  10.225 0.700 10.385 2.560 ;
        RECT  10.115 0.700 10.225 0.960 ;
        RECT  9.365 2.400 10.225 2.560 ;
        RECT  9.205 0.700 9.365 2.560 ;
        RECT  9.095 0.700 9.205 0.960 ;
        RECT  6.250 2.400 9.205 2.560 ;
        RECT  8.235 1.690 8.395 1.850 ;
        RECT  8.075 0.375 8.235 1.850 ;
        RECT  7.210 0.375 8.075 0.535 ;
        RECT  7.210 1.690 7.370 1.850 ;
        RECT  7.050 0.375 7.210 1.850 ;
        RECT  6.315 0.375 7.050 0.535 ;
        RECT  6.350 1.230 6.500 1.490 ;
        RECT  6.310 1.230 6.350 1.905 ;
        RECT  6.155 0.375 6.315 0.590 ;
        RECT  6.150 0.770 6.310 1.905 ;
        RECT  6.090 2.085 6.250 2.560 ;
        RECT  4.785 0.430 6.155 0.590 ;
        RECT  4.900 0.770 6.150 0.930 ;
        RECT  5.010 1.745 6.150 1.905 ;
        RECT  4.180 2.085 6.090 2.245 ;
        RECT  4.625 0.430 4.785 0.630 ;
        RECT  3.560 0.470 4.625 0.630 ;
        RECT  4.020 0.810 4.180 2.340 ;
        RECT  3.920 0.810 4.020 0.970 ;
        RECT  3.920 1.740 4.020 2.340 ;
        RECT  3.100 1.740 3.920 1.900 ;
        RECT  3.560 1.225 3.780 1.485 ;
        RECT  3.400 0.470 3.560 1.485 ;
        RECT  2.475 0.470 3.400 0.630 ;
        RECT  3.180 1.225 3.400 1.485 ;
        RECT  3.000 0.810 3.100 0.970 ;
        RECT  3.000 1.740 3.100 2.340 ;
        RECT  2.840 0.810 3.000 2.340 ;
        RECT  2.315 0.470 2.475 1.920 ;
        RECT  2.020 0.830 2.315 0.990 ;
        RECT  2.020 1.760 2.315 1.920 ;
        RECT  1.760 0.390 2.020 0.990 ;
        RECT  1.760 1.760 2.020 2.435 ;
        RECT  0.940 0.830 1.760 0.990 ;
        RECT  0.940 1.760 1.760 1.920 ;
        RECT  0.680 0.375 0.940 0.990 ;
        RECT  0.680 1.760 0.940 2.440 ;
    END
END XOR2X8MTH

MACRO XOR2XLMTH
    CLASS CORE ;
    FOREIGN XOR2XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.100 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.445 1.290 3.590 1.945 ;
        RECT  3.285 0.765 3.445 1.945 ;
        RECT  3.185 0.765 3.285 1.025 ;
        END
        AntennaDiffArea 0.238 ;
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.205 0.585 1.580 ;
        END
        AntennaGateArea 0.0702 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  1.585 1.215 1.950 1.830 ;
        END
        AntennaGateArea 0.1066 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.715 -0.130 4.100 0.130 ;
        RECT  0.775 -0.130 1.715 0.280 ;
        RECT  0.000 -0.130 0.775 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  1.750 2.740 4.100 3.000 ;
        RECT  0.810 2.465 1.750 3.000 ;
        RECT  0.000 2.740 0.810 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  3.815 0.335 3.975 2.515 ;
        RECT  3.715 0.335 3.815 0.595 ;
        RECT  3.715 2.125 3.815 2.515 ;
        RECT  1.405 2.125 3.715 2.285 ;
        RECT  2.795 0.475 2.955 1.945 ;
        RECT  2.625 0.475 2.795 1.025 ;
        RECT  2.695 1.685 2.795 1.945 ;
        RECT  0.935 0.475 2.625 0.635 ;
        RECT  2.445 1.245 2.570 1.505 ;
        RECT  2.285 0.815 2.445 1.920 ;
        RECT  2.105 0.815 2.285 0.975 ;
        RECT  2.185 1.760 2.285 1.920 ;
        RECT  1.245 0.815 1.405 2.285 ;
        RECT  1.145 0.815 1.245 0.975 ;
        RECT  1.195 1.685 1.245 1.945 ;
        RECT  0.935 1.225 1.015 1.485 ;
        RECT  0.775 0.475 0.935 1.920 ;
        RECT  0.385 0.865 0.775 1.025 ;
        RECT  0.125 1.760 0.775 1.920 ;
        RECT  0.125 0.765 0.385 1.025 ;
    END
END XOR2XLMTH

MACRO XOR3X1MTH
    CLASS CORE ;
    FOREIGN XOR3X1MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.950 0.755 8.110 2.005 ;
        RECT  7.815 0.755 7.950 1.015 ;
        RECT  7.815 1.700 7.950 2.005 ;
        END
        AntennaDiffArea 0.333 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.570 2.110 7.060 2.490 ;
        END
        AntennaGateArea 0.1937 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.120 4.820 1.740 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.555 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.880 -0.130 8.200 0.130 ;
        RECT  7.280 -0.130 7.880 0.250 ;
        RECT  4.840 -0.130 7.280 0.130 ;
        RECT  4.580 -0.130 4.840 0.860 ;
        RECT  2.810 -0.130 4.580 0.130 ;
        RECT  2.650 -0.130 2.810 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.995 2.740 8.200 3.000 ;
        RECT  7.395 2.555 7.995 3.000 ;
        RECT  4.820 2.740 7.395 3.000 ;
        RECT  4.600 2.265 4.820 3.000 ;
        RECT  2.545 2.740 4.600 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.840 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.635 1.235 7.765 1.495 ;
        RECT  7.475 0.430 7.635 1.495 ;
        RECT  7.035 0.430 7.475 0.590 ;
        RECT  7.025 1.735 7.085 1.895 ;
        RECT  6.875 0.310 7.035 0.590 ;
        RECT  6.755 0.815 7.025 1.895 ;
        RECT  5.900 0.310 6.875 0.470 ;
        RECT  6.710 0.815 6.755 0.975 ;
        RECT  6.535 1.245 6.755 1.505 ;
        RECT  6.355 1.735 6.575 1.895 ;
        RECT  6.355 0.655 6.460 0.925 ;
        RECT  6.195 0.655 6.355 2.560 ;
        RECT  5.160 2.400 6.195 2.560 ;
        RECT  5.900 1.825 6.015 2.085 ;
        RECT  5.740 0.310 5.900 2.085 ;
        RECT  5.400 0.645 5.560 2.080 ;
        RECT  5.180 0.645 5.400 0.905 ;
        RECT  5.340 1.820 5.400 2.080 ;
        RECT  5.160 1.265 5.220 1.525 ;
        RECT  5.000 1.265 5.160 2.560 ;
        RECT  4.420 1.925 5.000 2.085 ;
        RECT  4.260 1.925 4.420 2.560 ;
        RECT  4.240 0.310 4.400 1.745 ;
        RECT  2.885 2.400 4.260 2.560 ;
        RECT  3.430 0.310 4.240 0.470 ;
        RECT  4.080 1.585 4.240 1.745 ;
        RECT  3.920 1.585 4.080 2.220 ;
        RECT  3.900 0.650 4.060 1.385 ;
        RECT  3.230 2.060 3.920 2.220 ;
        RECT  3.740 1.225 3.900 1.385 ;
        RECT  3.580 1.225 3.740 1.880 ;
        RECT  2.470 0.885 3.720 1.045 ;
        RECT  1.875 1.225 3.580 1.385 ;
        RECT  3.170 0.310 3.430 0.675 ;
        RECT  3.070 1.565 3.230 2.220 ;
        RECT  1.865 1.565 3.070 1.725 ;
        RECT  2.725 1.905 2.885 2.560 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.895 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.675 2.130 0.935 ;
        RECT  1.405 2.320 2.045 2.480 ;
        RECT  1.695 0.775 1.970 0.935 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.355 2.095 1.405 2.480 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  1.145 2.095 1.195 2.355 ;
        RECT  0.735 0.310 0.895 2.410 ;
        RECT  0.635 0.460 0.735 0.720 ;
        RECT  0.635 1.810 0.735 2.410 ;
    END
END XOR3X1MTH

MACRO XOR3X2MTH
    CLASS CORE ;
    FOREIGN XOR3X2MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.200 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.945 0.415 8.105 2.405 ;
        RECT  7.815 0.415 7.945 1.015 ;
        RECT  7.815 1.805 7.945 2.405 ;
        END
        AntennaDiffArea 0.537 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  6.625 2.110 7.000 2.530 ;
        END
        AntennaGateArea 0.2457 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.120 4.820 1.705 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.505 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 -0.130 8.200 0.130 ;
        RECT  7.275 -0.130 7.535 0.250 ;
        RECT  4.840 -0.130 7.275 0.130 ;
        RECT  4.580 -0.130 4.840 0.840 ;
        RECT  2.810 -0.130 4.580 0.130 ;
        RECT  2.650 -0.130 2.810 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.535 2.740 8.200 3.000 ;
        RECT  7.275 2.265 7.535 3.000 ;
        RECT  4.820 2.740 7.275 3.000 ;
        RECT  4.660 2.265 4.820 3.000 ;
        RECT  2.545 2.740 4.660 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  7.635 1.235 7.765 1.495 ;
        RECT  7.475 0.430 7.635 1.495 ;
        RECT  7.095 0.430 7.475 0.590 ;
        RECT  6.935 0.310 7.095 0.590 ;
        RECT  7.045 1.735 7.085 1.895 ;
        RECT  6.755 0.815 7.045 1.895 ;
        RECT  5.900 0.310 6.935 0.470 ;
        RECT  6.710 0.815 6.755 0.975 ;
        RECT  6.535 1.245 6.755 1.505 ;
        RECT  6.355 1.735 6.575 1.895 ;
        RECT  6.355 0.650 6.460 0.810 ;
        RECT  6.195 0.650 6.355 2.560 ;
        RECT  5.160 2.400 6.195 2.560 ;
        RECT  5.900 1.905 6.015 2.165 ;
        RECT  5.740 0.310 5.900 2.165 ;
        RECT  5.400 0.525 5.560 2.220 ;
        RECT  5.180 0.525 5.400 0.785 ;
        RECT  5.340 1.960 5.400 2.220 ;
        RECT  5.160 1.265 5.220 1.525 ;
        RECT  5.000 1.265 5.160 2.560 ;
        RECT  4.480 1.925 5.000 2.085 ;
        RECT  4.320 1.925 4.480 2.560 ;
        RECT  4.240 0.310 4.400 1.745 ;
        RECT  2.885 2.400 4.320 2.560 ;
        RECT  3.430 0.310 4.240 0.470 ;
        RECT  4.140 1.585 4.240 1.745 ;
        RECT  3.980 1.585 4.140 2.220 ;
        RECT  3.900 0.655 4.060 1.385 ;
        RECT  3.290 2.060 3.980 2.220 ;
        RECT  3.800 1.225 3.900 1.385 ;
        RECT  3.640 1.225 3.800 1.880 ;
        RECT  2.470 0.885 3.720 1.045 ;
        RECT  1.875 1.225 3.640 1.385 ;
        RECT  3.170 0.310 3.430 0.675 ;
        RECT  3.130 1.565 3.290 2.220 ;
        RECT  1.865 1.565 3.130 1.725 ;
        RECT  2.725 1.905 2.885 2.560 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.845 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.675 2.130 0.935 ;
        RECT  1.405 2.320 2.045 2.480 ;
        RECT  1.695 0.775 1.970 0.935 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.775 1.695 1.725 ;
        RECT  1.300 1.865 1.405 2.480 ;
        RECT  1.300 0.650 1.355 0.910 ;
        RECT  1.140 0.650 1.300 2.480 ;
        RECT  0.845 1.860 0.895 2.460 ;
        RECT  0.685 0.310 0.845 2.460 ;
        RECT  0.635 1.860 0.685 2.460 ;
    END
END XOR3X2MTH

MACRO XOR3X4MTH
    CLASS CORE ;
    FOREIGN XOR3X4MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.430 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  8.685 0.380 8.865 2.410 ;
        RECT  8.535 0.380 8.685 0.980 ;
        RECT  8.535 1.680 8.685 2.410 ;
        RECT  8.260 1.680 8.535 1.950 ;
        END
        AntennaDiffArea 0.6 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.280 2.075 7.815 2.495 ;
        END
        AntennaGateArea 0.247 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.580 1.070 4.820 1.690 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.555 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 -0.130 9.430 0.130 ;
        RECT  9.045 -0.130 9.305 0.990 ;
        RECT  8.255 -0.130 9.045 0.130 ;
        RECT  7.995 -0.130 8.255 0.295 ;
        RECT  5.675 -0.130 7.995 0.130 ;
        RECT  5.415 -0.130 5.675 0.565 ;
        RECT  2.810 -0.130 5.415 0.130 ;
        RECT  2.650 -0.130 2.810 0.705 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.955 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  9.305 2.740 9.430 3.000 ;
        RECT  9.045 1.790 9.305 3.000 ;
        RECT  8.255 2.740 9.045 3.000 ;
        RECT  7.995 2.130 8.255 3.000 ;
        RECT  5.610 2.740 7.995 3.000 ;
        RECT  5.350 2.585 5.610 3.000 ;
        RECT  2.545 2.740 5.350 3.000 ;
        RECT  2.385 2.245 2.545 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.815 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.355 1.235 8.505 1.495 ;
        RECT  8.195 0.475 8.355 1.495 ;
        RECT  7.815 0.475 8.195 0.635 ;
        RECT  7.655 0.310 7.815 0.635 ;
        RECT  7.565 0.815 7.725 1.895 ;
        RECT  6.645 0.310 7.655 0.470 ;
        RECT  7.455 0.815 7.565 0.975 ;
        RECT  7.290 1.315 7.565 1.475 ;
        RECT  7.420 1.735 7.565 1.895 ;
        RECT  7.130 1.315 7.290 1.575 ;
        RECT  7.055 0.655 7.205 0.815 ;
        RECT  6.950 1.765 7.170 1.925 ;
        RECT  6.950 0.655 7.055 1.110 ;
        RECT  6.895 0.655 6.950 2.405 ;
        RECT  6.790 0.950 6.895 2.405 ;
        RECT  5.760 2.245 6.790 2.405 ;
        RECT  6.610 0.310 6.645 0.840 ;
        RECT  6.450 0.310 6.610 2.065 ;
        RECT  6.100 0.505 6.185 0.915 ;
        RECT  5.940 0.505 6.100 2.065 ;
        RECT  5.925 0.505 5.940 0.915 ;
        RECT  5.165 0.755 5.925 0.915 ;
        RECT  5.600 1.265 5.760 2.405 ;
        RECT  5.380 1.265 5.600 1.525 ;
        RECT  4.470 2.220 5.600 2.380 ;
        RECT  5.160 0.505 5.165 0.915 ;
        RECT  5.000 0.505 5.160 2.035 ;
        RECT  4.905 0.505 5.000 0.765 ;
        RECT  4.810 1.875 5.000 2.035 ;
        RECT  4.310 2.220 4.470 2.510 ;
        RECT  4.240 0.310 4.400 1.745 ;
        RECT  2.885 2.350 4.310 2.510 ;
        RECT  3.430 0.310 4.240 0.470 ;
        RECT  4.130 1.585 4.240 1.745 ;
        RECT  3.970 1.585 4.130 2.170 ;
        RECT  3.900 0.650 4.060 1.385 ;
        RECT  3.230 2.010 3.970 2.170 ;
        RECT  3.790 1.225 3.900 1.385 ;
        RECT  3.630 1.225 3.790 1.830 ;
        RECT  2.470 0.885 3.720 1.045 ;
        RECT  1.875 1.225 3.630 1.385 ;
        RECT  3.530 1.670 3.630 1.830 ;
        RECT  3.170 0.310 3.430 0.675 ;
        RECT  3.070 1.565 3.230 2.170 ;
        RECT  1.865 1.565 3.070 1.725 ;
        RECT  2.725 1.905 2.885 2.510 ;
        RECT  2.205 1.905 2.725 2.065 ;
        RECT  2.310 0.310 2.470 1.045 ;
        RECT  0.895 0.310 2.310 0.470 ;
        RECT  2.045 1.905 2.205 2.480 ;
        RECT  1.970 0.705 2.130 0.965 ;
        RECT  1.355 2.320 2.045 2.480 ;
        RECT  1.695 0.805 1.970 0.965 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.805 1.695 1.725 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  0.735 0.310 0.895 2.455 ;
        RECT  0.635 0.520 0.735 0.780 ;
        RECT  0.635 1.855 0.735 2.455 ;
    END
END XOR3X4MTH

MACRO XOR3X8MTH
    CLASS CORE ;
    FOREIGN XOR3X8MTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.070 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  10.145 0.415 10.465 2.370 ;
        RECT  9.480 1.235 10.145 1.585 ;
        RECT  9.250 0.415 9.480 2.390 ;
        RECT  9.155 0.415 9.250 1.015 ;
        RECT  9.155 1.790 9.250 2.390 ;
        END
        AntennaDiffArea 1.2 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.985 2.075 8.510 2.400 ;
        END
        AntennaGateArea 0.247 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  4.345 1.175 4.820 1.610 ;
        END
        AntennaGateArea 0.247 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.040 0.355 1.580 ;
        END
        AntennaGateArea 0.2054 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 -0.130 11.070 0.130 ;
        RECT  10.685 -0.130 10.945 0.990 ;
        RECT  9.925 -0.130 10.685 0.130 ;
        RECT  9.665 -0.130 9.925 0.955 ;
        RECT  8.875 -0.130 9.665 0.130 ;
        RECT  8.615 -0.130 8.875 0.250 ;
        RECT  6.345 -0.130 8.615 0.130 ;
        RECT  6.085 -0.130 6.345 0.565 ;
        RECT  5.325 -0.130 6.085 0.130 ;
        RECT  5.065 -0.130 5.325 0.565 ;
        RECT  2.655 -0.130 5.065 0.130 ;
        RECT  2.495 -0.130 2.655 0.705 ;
        RECT  0.000 -0.130 2.495 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  10.945 2.740 11.070 3.000 ;
        RECT  10.685 1.805 10.945 3.000 ;
        RECT  9.925 2.740 10.685 3.000 ;
        RECT  9.665 1.915 9.925 3.000 ;
        RECT  8.875 2.740 9.665 3.000 ;
        RECT  8.615 2.550 8.875 3.000 ;
        RECT  6.315 2.740 8.615 3.000 ;
        RECT  6.055 2.530 6.315 3.000 ;
        RECT  5.235 2.740 6.055 3.000 ;
        RECT  4.975 2.530 5.235 3.000 ;
        RECT  2.435 2.740 4.975 3.000 ;
        RECT  2.275 2.245 2.435 3.000 ;
        RECT  0.000 2.740 2.275 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  8.975 1.235 9.070 1.495 ;
        RECT  8.815 0.430 8.975 1.495 ;
        RECT  8.385 0.430 8.815 0.590 ;
        RECT  8.385 0.815 8.440 0.975 ;
        RECT  8.225 0.310 8.385 0.590 ;
        RECT  8.125 0.815 8.385 1.895 ;
        RECT  7.370 0.310 8.225 0.470 ;
        RECT  7.955 1.315 8.125 1.575 ;
        RECT  7.775 0.650 7.930 0.865 ;
        RECT  7.775 1.740 7.875 1.930 ;
        RECT  7.615 0.650 7.775 2.350 ;
        RECT  6.320 2.190 7.615 2.350 ;
        RECT  7.210 0.310 7.370 2.010 ;
        RECT  7.105 1.850 7.210 2.010 ;
        RECT  6.755 0.495 6.910 0.910 ;
        RECT  6.755 1.850 6.855 2.010 ;
        RECT  6.595 0.495 6.755 2.010 ;
        RECT  5.835 0.750 6.595 0.910 ;
        RECT  6.320 1.265 6.415 1.525 ;
        RECT  6.160 1.265 6.320 2.350 ;
        RECT  5.475 1.265 6.160 1.525 ;
        RECT  4.305 2.190 6.160 2.350 ;
        RECT  5.575 0.495 5.835 0.910 ;
        RECT  5.270 1.850 5.775 2.010 ;
        RECT  5.270 0.750 5.575 0.910 ;
        RECT  5.110 0.750 5.270 2.010 ;
        RECT  4.815 0.750 5.110 0.910 ;
        RECT  4.435 1.850 5.110 2.010 ;
        RECT  4.555 0.495 4.815 0.910 ;
        RECT  4.145 2.190 4.305 2.560 ;
        RECT  4.005 0.310 4.165 1.745 ;
        RECT  2.775 2.400 4.145 2.560 ;
        RECT  3.275 0.310 4.005 0.470 ;
        RECT  3.965 1.585 4.005 1.745 ;
        RECT  3.805 1.585 3.965 2.220 ;
        RECT  3.665 0.650 3.825 1.385 ;
        RECT  3.115 2.060 3.805 2.220 ;
        RECT  3.625 1.225 3.665 1.385 ;
        RECT  3.465 1.225 3.625 1.880 ;
        RECT  1.765 1.225 3.465 1.385 ;
        RECT  3.295 0.785 3.455 1.045 ;
        RECT  2.315 0.885 3.295 1.045 ;
        RECT  3.015 0.310 3.275 0.605 ;
        RECT  2.955 1.565 3.115 2.220 ;
        RECT  1.755 1.565 2.955 1.725 ;
        RECT  2.615 1.905 2.775 2.560 ;
        RECT  2.095 1.905 2.615 2.065 ;
        RECT  2.155 0.310 2.315 1.045 ;
        RECT  0.735 0.310 2.155 0.470 ;
        RECT  1.935 1.905 2.095 2.480 ;
        RECT  1.815 0.675 1.975 0.935 ;
        RECT  1.245 2.320 1.935 2.480 ;
        RECT  1.585 0.775 1.815 0.935 ;
        RECT  1.595 1.565 1.755 2.140 ;
        RECT  1.585 1.565 1.595 1.725 ;
        RECT  1.425 0.775 1.585 1.725 ;
        RECT  1.085 0.650 1.245 2.480 ;
        RECT  0.735 1.810 0.785 2.410 ;
        RECT  0.575 0.310 0.735 2.410 ;
        RECT  0.525 1.810 0.575 2.410 ;
    END
END XOR3X8MTH

MACRO XOR3XLMTH
    CLASS CORE ;
    FOREIGN XOR3XLMTH 0.000 0.000  ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.380 BY 2.870 ;
    SYMMETRY X Y ;
    SITE TSM130NMMETROSITE ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER METAL1 ;
        RECT  7.120 0.765 7.280 1.990 ;
        RECT  6.995 0.765 7.120 1.025 ;
        RECT  6.995 1.700 7.120 1.990 ;
        END
        AntennaDiffArea 0.236 ;
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  5.780 2.110 6.240 2.490 ;
        END
        AntennaGateArea 0.1586 ;
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  3.570 1.120 4.000 1.635 ;
        END
        AntennaGateArea 0.1794 ;
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER METAL1 ;
        RECT  0.100 1.170 0.555 1.580 ;
        END
        AntennaGateArea 0.1378 ;
    END A
    PIN VSS
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.090 -0.130 7.380 0.130 ;
        RECT  6.490 -0.130 7.090 0.285 ;
        RECT  4.670 -0.130 6.490 0.130 ;
        RECT  3.990 -0.130 4.670 0.330 ;
        RECT  3.730 -0.130 3.990 0.910 ;
        RECT  2.910 -0.130 3.730 0.130 ;
        RECT  2.650 -0.130 2.910 0.655 ;
        RECT  0.385 -0.130 2.650 0.130 ;
        RECT  0.125 -0.130 0.385 0.825 ;
        RECT  0.000 -0.130 0.125 0.130 ;
        END
    END VSS
    PIN VDD
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER METAL1 ;
        RECT  7.090 2.740 7.380 3.000 ;
        RECT  6.490 2.315 7.090 3.000 ;
        RECT  3.950 2.740 6.490 3.000 ;
        RECT  3.690 2.490 3.950 3.000 ;
        RECT  2.645 2.740 3.690 3.000 ;
        RECT  2.385 2.085 2.645 3.000 ;
        RECT  0.385 2.740 2.385 3.000 ;
        RECT  0.125 1.895 0.385 3.000 ;
        RECT  0.000 2.740 0.125 3.000 ;
        END
    END VDD
    OBS
        LAYER METAL1 ;
        RECT  6.815 1.235 6.885 1.495 ;
        RECT  6.655 0.475 6.815 1.495 ;
        RECT  6.130 0.475 6.655 0.635 ;
        RECT  6.625 1.235 6.655 1.495 ;
        RECT  5.920 0.815 6.190 1.895 ;
        RECT  5.970 0.310 6.130 0.635 ;
        RECT  5.110 0.310 5.970 0.470 ;
        RECT  5.630 1.310 5.920 1.570 ;
        RECT  5.450 0.650 5.670 0.910 ;
        RECT  5.450 1.765 5.620 2.025 ;
        RECT  5.290 0.650 5.450 2.560 ;
        RECT  4.390 2.400 5.290 2.560 ;
        RECT  4.950 0.310 5.110 2.060 ;
        RECT  4.430 0.650 4.590 1.945 ;
        RECT  4.330 0.650 4.430 0.910 ;
        RECT  4.330 1.685 4.430 1.945 ;
        RECT  4.130 2.150 4.390 2.560 ;
        RECT  2.990 2.150 4.130 2.310 ;
        RECT  3.330 0.650 3.390 1.565 ;
        RECT  3.230 0.650 3.330 1.945 ;
        RECT  3.190 0.650 3.230 0.910 ;
        RECT  3.170 1.405 3.230 1.945 ;
        RECT  2.205 1.405 3.170 1.565 ;
        RECT  2.950 1.065 3.050 1.225 ;
        RECT  2.830 1.745 2.990 2.310 ;
        RECT  2.790 0.835 2.950 1.225 ;
        RECT  2.205 1.745 2.830 1.905 ;
        RECT  2.470 0.835 2.790 0.995 ;
        RECT  2.310 0.310 2.470 0.995 ;
        RECT  0.895 0.310 2.310 0.470 ;
        RECT  2.045 1.145 2.205 1.565 ;
        RECT  2.045 1.745 2.205 2.480 ;
        RECT  1.970 0.690 2.130 0.950 ;
        RECT  1.875 1.145 2.045 1.305 ;
        RECT  1.355 2.320 2.045 2.480 ;
        RECT  1.695 0.790 1.970 0.950 ;
        RECT  1.705 1.565 1.865 2.140 ;
        RECT  1.695 1.565 1.705 1.725 ;
        RECT  1.535 0.790 1.695 1.725 ;
        RECT  1.195 0.650 1.355 2.480 ;
        RECT  0.735 0.310 0.895 2.155 ;
        RECT  0.635 0.560 0.735 0.820 ;
        RECT  0.635 1.895 0.735 2.155 ;
    END
END XOR3XLMTH

END LIBRARY
